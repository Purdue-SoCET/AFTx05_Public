`include "memory_blocks_if.vh"

module SOC_ROM(memory_blocks_if.rom blkif);

parameter ROM_TOP = 16'h2000;
parameter ROM_BOTTOM  = 16'h3b;

logic [31:0] addr;

assign addr = blkif.addr >> 2; // ROM is byte addressed

assign blkif.rom_active = addr >= ROM_BOTTOM && addr < ROM_TOP;
assign blkif.rom_wait = 1'b0;

always_comb begin
        case (addr)
          16'h0080 : blkif.rom_rdata <= 32'h23200000;
          16'h0081 : blkif.rom_rdata <= 32'hb7000080;
          16'h0082 : blkif.rom_rdata <= 32'h93808000;
          16'h0083 : blkif.rom_rdata <= 32'h23a00000;
          16'h0084 : blkif.rom_rdata <= 32'hb7000080;
          16'h0085 : blkif.rom_rdata <= 32'h93804000;
          16'h0086 : blkif.rom_rdata <= 32'h13000000;
          16'h0087 : blkif.rom_rdata <= 32'h13000000;
          16'h0088 : blkif.rom_rdata <= 32'h13000000;
          16'h0089 : blkif.rom_rdata <= 32'h13000000;
          16'h008a : blkif.rom_rdata <= 32'h13000000;
          16'h008b : blkif.rom_rdata <= 32'h13000000;
          16'h008c : blkif.rom_rdata <= 32'h13000000;
          16'h008d : blkif.rom_rdata <= 32'h13000000;
          16'h008e : blkif.rom_rdata <= 32'h03a10000;
          16'h008f : blkif.rom_rdata <= 32'h13711100;
          16'h0090 : blkif.rom_rdata <= 32'h63100102;
          16'h0091 : blkif.rom_rdata <= 32'h83210000;
          16'h0092 : blkif.rom_rdata <= 32'he38801fe;
          16'h0093 : blkif.rom_rdata <= 32'hb7000080;
          16'h0094 : blkif.rom_rdata <= 32'h93808000;
          16'h0095 : blkif.rom_rdata <= 32'h1301f00f;
          16'h0096 : blkif.rom_rdata <= 32'h23a02000;
          16'h0097 : blkif.rom_rdata <= 32'h67820100;
          16'h0098 : blkif.rom_rdata <= 32'hb7000080;
          16'h0099 : blkif.rom_rdata <= 32'h93808000;
          16'h009a : blkif.rom_rdata <= 32'h1301f00f;
          16'h009b : blkif.rom_rdata <= 32'h23a02000;
          16'h009c : blkif.rom_rdata <= 32'hb7000080;
          16'h009d : blkif.rom_rdata <= 32'h93804000;
          16'h009e : blkif.rom_rdata <= 32'h13012000;
          16'h009f : blkif.rom_rdata <= 32'h23a02000;
          16'h00a0 : blkif.rom_rdata <= 32'h93000000;
          16'h00a1 : blkif.rom_rdata <= 32'h13010000;
          16'h00a2 : blkif.rom_rdata <= 32'hb3812000;
          16'h00a3 : blkif.rom_rdata <= 32'h930e0000;
          16'h00a4 : blkif.rom_rdata <= 32'h130e2000;
          16'h00a5 : blkif.rom_rdata <= 32'h6384d101;
          16'h00a6 : blkif.rom_rdata <= 32'h6f50404d;
          16'h00a7 : blkif.rom_rdata <= 32'hb7000080;
          16'h00a8 : blkif.rom_rdata <= 32'h93804000;
          16'h00a9 : blkif.rom_rdata <= 32'h13013000;
          16'h00aa : blkif.rom_rdata <= 32'h23a02000;
          16'h00ab : blkif.rom_rdata <= 32'h9300f0ff;
          16'h00ac : blkif.rom_rdata <= 32'h1301f0ff;
          16'h00ad : blkif.rom_rdata <= 32'hb3812000;
          16'h00ae : blkif.rom_rdata <= 32'h930ee0ff;
          16'h00af : blkif.rom_rdata <= 32'h130e3000;
          16'h00b0 : blkif.rom_rdata <= 32'h6384d101;
          16'h00b1 : blkif.rom_rdata <= 32'h6f50804a;
          16'h00b2 : blkif.rom_rdata <= 32'hb7000080;
          16'h00b3 : blkif.rom_rdata <= 32'h93804000;
          16'h00b4 : blkif.rom_rdata <= 32'h13010001;
          16'h00b5 : blkif.rom_rdata <= 32'h23a02000;
          16'h00b6 : blkif.rom_rdata <= 32'h93001000;
          16'h00b7 : blkif.rom_rdata <= 32'h37010080;
          16'h00b8 : blkif.rom_rdata <= 32'h1301f1ff;
          16'h00b9 : blkif.rom_rdata <= 32'hb3812000;
          16'h00ba : blkif.rom_rdata <= 32'hb70e0080;
          16'h00bb : blkif.rom_rdata <= 32'h130e0001;
          16'h00bc : blkif.rom_rdata <= 32'h6384d101;
          16'h00bd : blkif.rom_rdata <= 32'h6f508047;
          16'h00be : blkif.rom_rdata <= 32'hb7000080;
          16'h00bf : blkif.rom_rdata <= 32'h93804000;
          16'h00c0 : blkif.rom_rdata <= 32'h13011001;
          16'h00c1 : blkif.rom_rdata <= 32'h23a02000;
          16'h00c2 : blkif.rom_rdata <= 32'h9300d000;
          16'h00c3 : blkif.rom_rdata <= 32'h1301b000;
          16'h00c4 : blkif.rom_rdata <= 32'hb3802000;
          16'h00c5 : blkif.rom_rdata <= 32'h930e8001;
          16'h00c6 : blkif.rom_rdata <= 32'h130e1001;
          16'h00c7 : blkif.rom_rdata <= 32'h6384d001;
          16'h00c8 : blkif.rom_rdata <= 32'h6f50c044;
          16'h00c9 : blkif.rom_rdata <= 32'hb7000080;
          16'h00ca : blkif.rom_rdata <= 32'h93804000;
          16'h00cb : blkif.rom_rdata <= 32'h13012001;
          16'h00cc : blkif.rom_rdata <= 32'h23a02000;
          16'h00cd : blkif.rom_rdata <= 32'h9300e000;
          16'h00ce : blkif.rom_rdata <= 32'h1301b000;
          16'h00cf : blkif.rom_rdata <= 32'h33812000;
          16'h00d0 : blkif.rom_rdata <= 32'h930e9001;
          16'h00d1 : blkif.rom_rdata <= 32'h130e2001;
          16'h00d2 : blkif.rom_rdata <= 32'h6304d101;
          16'h00d3 : blkif.rom_rdata <= 32'h6f500042;
          16'h00d4 : blkif.rom_rdata <= 32'hb7000080;
          16'h00d5 : blkif.rom_rdata <= 32'h93804000;
          16'h00d6 : blkif.rom_rdata <= 32'h13013001;
          16'h00d7 : blkif.rom_rdata <= 32'h23a02000;
          16'h00d8 : blkif.rom_rdata <= 32'h9300d000;
          16'h00d9 : blkif.rom_rdata <= 32'hb3801000;
          16'h00da : blkif.rom_rdata <= 32'h930ea001;
          16'h00db : blkif.rom_rdata <= 32'h130e3001;
          16'h00dc : blkif.rom_rdata <= 32'h6384d001;
          16'h00dd : blkif.rom_rdata <= 32'h6f50803f;
          16'h00de : blkif.rom_rdata <= 32'hb7000080;
          16'h00df : blkif.rom_rdata <= 32'h93804000;
          16'h00e0 : blkif.rom_rdata <= 32'h13014001;
          16'h00e1 : blkif.rom_rdata <= 32'h23a02000;
          16'h00e2 : blkif.rom_rdata <= 32'h13020000;
          16'h00e3 : blkif.rom_rdata <= 32'h9300d000;
          16'h00e4 : blkif.rom_rdata <= 32'h1301b000;
          16'h00e5 : blkif.rom_rdata <= 32'hb3812000;
          16'h00e6 : blkif.rom_rdata <= 32'h13830100;
          16'h00e7 : blkif.rom_rdata <= 32'h13021200;
          16'h00e8 : blkif.rom_rdata <= 32'h93022000;
          16'h00e9 : blkif.rom_rdata <= 32'he31452fe;
          16'h00ea : blkif.rom_rdata <= 32'h930e8001;
          16'h00eb : blkif.rom_rdata <= 32'h130e4001;
          16'h00ec : blkif.rom_rdata <= 32'h6304d301;
          16'h00ed : blkif.rom_rdata <= 32'h6f50803b;
          16'h00ee : blkif.rom_rdata <= 32'hb7000080;
          16'h00ef : blkif.rom_rdata <= 32'h93804000;
          16'h00f0 : blkif.rom_rdata <= 32'h13016001;
          16'h00f1 : blkif.rom_rdata <= 32'h23a02000;
          16'h00f2 : blkif.rom_rdata <= 32'h13020000;
          16'h00f3 : blkif.rom_rdata <= 32'h9300f000;
          16'h00f4 : blkif.rom_rdata <= 32'h1301b000;
          16'h00f5 : blkif.rom_rdata <= 32'hb3812000;
          16'h00f6 : blkif.rom_rdata <= 32'h13000000;
          16'h00f7 : blkif.rom_rdata <= 32'h13000000;
          16'h00f8 : blkif.rom_rdata <= 32'h13830100;
          16'h00f9 : blkif.rom_rdata <= 32'h13021200;
          16'h00fa : blkif.rom_rdata <= 32'h93022000;
          16'h00fb : blkif.rom_rdata <= 32'he31052fe;
          16'h00fc : blkif.rom_rdata <= 32'h930ea001;
          16'h00fd : blkif.rom_rdata <= 32'h130e6001;
          16'h00fe : blkif.rom_rdata <= 32'h6304d301;
          16'h00ff : blkif.rom_rdata <= 32'h6f500037;
          16'h0100 : blkif.rom_rdata <= 32'hb7000080;
          16'h0101 : blkif.rom_rdata <= 32'h93804000;
          16'h0102 : blkif.rom_rdata <= 32'h13017001;
          16'h0103 : blkif.rom_rdata <= 32'h23a02000;
          16'h0104 : blkif.rom_rdata <= 32'h13020000;
          16'h0105 : blkif.rom_rdata <= 32'h9300d000;
          16'h0106 : blkif.rom_rdata <= 32'h1301b000;
          16'h0107 : blkif.rom_rdata <= 32'hb3812000;
          16'h0108 : blkif.rom_rdata <= 32'h13021200;
          16'h0109 : blkif.rom_rdata <= 32'h93022000;
          16'h010a : blkif.rom_rdata <= 32'he31652fe;
          16'h010b : blkif.rom_rdata <= 32'h930e8001;
          16'h010c : blkif.rom_rdata <= 32'h130e7001;
          16'h010d : blkif.rom_rdata <= 32'h6384d101;
          16'h010e : blkif.rom_rdata <= 32'h6f504033;
          16'h010f : blkif.rom_rdata <= 32'hb7000080;
          16'h0110 : blkif.rom_rdata <= 32'h93804000;
          16'h0111 : blkif.rom_rdata <= 32'h13018001;
          16'h0112 : blkif.rom_rdata <= 32'h23a02000;
          16'h0113 : blkif.rom_rdata <= 32'h13020000;
          16'h0114 : blkif.rom_rdata <= 32'h9300e000;
          16'h0115 : blkif.rom_rdata <= 32'h1301b000;
          16'h0116 : blkif.rom_rdata <= 32'h13000000;
          16'h0117 : blkif.rom_rdata <= 32'hb3812000;
          16'h0118 : blkif.rom_rdata <= 32'h13021200;
          16'h0119 : blkif.rom_rdata <= 32'h93022000;
          16'h011a : blkif.rom_rdata <= 32'he31452fe;
          16'h011b : blkif.rom_rdata <= 32'h930e9001;
          16'h011c : blkif.rom_rdata <= 32'h130e8001;
          16'h011d : blkif.rom_rdata <= 32'h6384d101;
          16'h011e : blkif.rom_rdata <= 32'h6f50402f;
          16'h011f : blkif.rom_rdata <= 32'hb7000080;
          16'h0120 : blkif.rom_rdata <= 32'h93804000;
          16'h0121 : blkif.rom_rdata <= 32'h1301c001;
          16'h0122 : blkif.rom_rdata <= 32'h23a02000;
          16'h0123 : blkif.rom_rdata <= 32'h13020000;
          16'h0124 : blkif.rom_rdata <= 32'h9300f000;
          16'h0125 : blkif.rom_rdata <= 32'h13000000;
          16'h0126 : blkif.rom_rdata <= 32'h13000000;
          16'h0127 : blkif.rom_rdata <= 32'h1301b000;
          16'h0128 : blkif.rom_rdata <= 32'hb3812000;
          16'h0129 : blkif.rom_rdata <= 32'h13021200;
          16'h012a : blkif.rom_rdata <= 32'h93022000;
          16'h012b : blkif.rom_rdata <= 32'he31252fe;
          16'h012c : blkif.rom_rdata <= 32'h930ea001;
          16'h012d : blkif.rom_rdata <= 32'h130ec001;
          16'h012e : blkif.rom_rdata <= 32'h6384d101;
          16'h012f : blkif.rom_rdata <= 32'h6f50002b;
          16'h0130 : blkif.rom_rdata <= 32'hb7000080;
          16'h0131 : blkif.rom_rdata <= 32'h93804000;
          16'h0132 : blkif.rom_rdata <= 32'h13012002;
          16'h0133 : blkif.rom_rdata <= 32'h23a02000;
          16'h0134 : blkif.rom_rdata <= 32'h13020000;
          16'h0135 : blkif.rom_rdata <= 32'h1301b000;
          16'h0136 : blkif.rom_rdata <= 32'h13000000;
          16'h0137 : blkif.rom_rdata <= 32'h13000000;
          16'h0138 : blkif.rom_rdata <= 32'h9300f000;
          16'h0139 : blkif.rom_rdata <= 32'hb3812000;
          16'h013a : blkif.rom_rdata <= 32'h13021200;
          16'h013b : blkif.rom_rdata <= 32'h93022000;
          16'h013c : blkif.rom_rdata <= 32'he31252fe;
          16'h013d : blkif.rom_rdata <= 32'h930ea001;
          16'h013e : blkif.rom_rdata <= 32'h130e2002;
          16'h013f : blkif.rom_rdata <= 32'h6384d101;
          16'h0140 : blkif.rom_rdata <= 32'h6f50c026;
          16'h0141 : blkif.rom_rdata <= 32'hb7000080;
          16'h0142 : blkif.rom_rdata <= 32'h93804000;
          16'h0143 : blkif.rom_rdata <= 32'h13013002;
          16'h0144 : blkif.rom_rdata <= 32'h23a02000;
          16'h0145 : blkif.rom_rdata <= 32'h9300f000;
          16'h0146 : blkif.rom_rdata <= 32'h33011000;
          16'h0147 : blkif.rom_rdata <= 32'h930ef000;
          16'h0148 : blkif.rom_rdata <= 32'h130e3002;
          16'h0149 : blkif.rom_rdata <= 32'h6304d101;
          16'h014a : blkif.rom_rdata <= 32'h6f504024;
          16'h014b : blkif.rom_rdata <= 32'hb7000080;
          16'h014c : blkif.rom_rdata <= 32'h93804000;
          16'h014d : blkif.rom_rdata <= 32'h13016002;
          16'h014e : blkif.rom_rdata <= 32'h23a02000;
          16'h014f : blkif.rom_rdata <= 32'h93000001;
          16'h0150 : blkif.rom_rdata <= 32'h1301e001;
          16'h0151 : blkif.rom_rdata <= 32'h33802000;
          16'h0152 : blkif.rom_rdata <= 32'h930e0000;
          16'h0153 : blkif.rom_rdata <= 32'h130e6002;
          16'h0154 : blkif.rom_rdata <= 32'h6304d001;
          16'h0155 : blkif.rom_rdata <= 32'h6f508021;
          16'h0156 : blkif.rom_rdata <= 32'hb7000080;
          16'h0157 : blkif.rom_rdata <= 32'h93804000;
          16'h0158 : blkif.rom_rdata <= 32'h13017002;
          16'h0159 : blkif.rom_rdata <= 32'h23a02000;
          16'h015a : blkif.rom_rdata <= 32'h93000000;
          16'h015b : blkif.rom_rdata <= 32'h93810000;
          16'h015c : blkif.rom_rdata <= 32'h930e0000;
          16'h015d : blkif.rom_rdata <= 32'h130e7002;
          16'h015e : blkif.rom_rdata <= 32'h6384d101;
          16'h015f : blkif.rom_rdata <= 32'h6f50001f;
          16'h0160 : blkif.rom_rdata <= 32'hb7000080;
          16'h0161 : blkif.rom_rdata <= 32'h93804000;
          16'h0162 : blkif.rom_rdata <= 32'h13019002;
          16'h0163 : blkif.rom_rdata <= 32'h23a02000;
          16'h0164 : blkif.rom_rdata <= 32'h93003000;
          16'h0165 : blkif.rom_rdata <= 32'h93817000;
          16'h0166 : blkif.rom_rdata <= 32'h930ea000;
          16'h0167 : blkif.rom_rdata <= 32'h130e9002;
          16'h0168 : blkif.rom_rdata <= 32'h6384d101;
          16'h0169 : blkif.rom_rdata <= 32'h6f50801c;
          16'h016a : blkif.rom_rdata <= 32'hb7000080;
          16'h016b : blkif.rom_rdata <= 32'h93804000;
          16'h016c : blkif.rom_rdata <= 32'h1301a002;
          16'h016d : blkif.rom_rdata <= 32'h23a02000;
          16'h016e : blkif.rom_rdata <= 32'h93000000;
          16'h016f : blkif.rom_rdata <= 32'h93810080;
          16'h0170 : blkif.rom_rdata <= 32'h930e0080;
          16'h0171 : blkif.rom_rdata <= 32'h130ea002;
          16'h0172 : blkif.rom_rdata <= 32'h6384d101;
          16'h0173 : blkif.rom_rdata <= 32'h6f50001a;
          16'h0174 : blkif.rom_rdata <= 32'hb7000080;
          16'h0175 : blkif.rom_rdata <= 32'h93804000;
          16'h0176 : blkif.rom_rdata <= 32'h1301c002;
          16'h0177 : blkif.rom_rdata <= 32'h23a02000;
          16'h0178 : blkif.rom_rdata <= 32'hb7000080;
          16'h0179 : blkif.rom_rdata <= 32'h93810080;
          16'h017a : blkif.rom_rdata <= 32'hb70e0080;
          16'h017b : blkif.rom_rdata <= 32'h938e0e80;
          16'h017c : blkif.rom_rdata <= 32'h130ec002;
          16'h017d : blkif.rom_rdata <= 32'h6384d101;
          16'h017e : blkif.rom_rdata <= 32'h6f504017;
          16'h017f : blkif.rom_rdata <= 32'hb7000080;
          16'h0180 : blkif.rom_rdata <= 32'h93804000;
          16'h0181 : blkif.rom_rdata <= 32'h13012003;
          16'h0182 : blkif.rom_rdata <= 32'h23a02000;
          16'h0183 : blkif.rom_rdata <= 32'h93000000;
          16'h0184 : blkif.rom_rdata <= 32'h9381f0ff;
          16'h0185 : blkif.rom_rdata <= 32'h930ef0ff;
          16'h0186 : blkif.rom_rdata <= 32'h130e2003;
          16'h0187 : blkif.rom_rdata <= 32'h6384d101;
          16'h0188 : blkif.rom_rdata <= 32'h6f50c014;
          16'h0189 : blkif.rom_rdata <= 32'hb7000080;
          16'h018a : blkif.rom_rdata <= 32'h93804000;
          16'h018b : blkif.rom_rdata <= 32'h13015003;
          16'h018c : blkif.rom_rdata <= 32'h23a02000;
          16'h018d : blkif.rom_rdata <= 32'hb7000080;
          16'h018e : blkif.rom_rdata <= 32'h9380f0ff;
          16'h018f : blkif.rom_rdata <= 32'h93811000;
          16'h0190 : blkif.rom_rdata <= 32'hb70e0080;
          16'h0191 : blkif.rom_rdata <= 32'h130e5003;
          16'h0192 : blkif.rom_rdata <= 32'h6384d101;
          16'h0193 : blkif.rom_rdata <= 32'h6f500012;
          16'h0194 : blkif.rom_rdata <= 32'hb7000080;
          16'h0195 : blkif.rom_rdata <= 32'h93804000;
          16'h0196 : blkif.rom_rdata <= 32'h13016003;
          16'h0197 : blkif.rom_rdata <= 32'h23a02000;
          16'h0198 : blkif.rom_rdata <= 32'h9300d000;
          16'h0199 : blkif.rom_rdata <= 32'h9380b000;
          16'h019a : blkif.rom_rdata <= 32'h930e8001;
          16'h019b : blkif.rom_rdata <= 32'h130e6003;
          16'h019c : blkif.rom_rdata <= 32'h6384d001;
          16'h019d : blkif.rom_rdata <= 32'h6f50800f;
          16'h019e : blkif.rom_rdata <= 32'hb7000080;
          16'h019f : blkif.rom_rdata <= 32'h93804000;
          16'h01a0 : blkif.rom_rdata <= 32'h13017003;
          16'h01a1 : blkif.rom_rdata <= 32'h23a02000;
          16'h01a2 : blkif.rom_rdata <= 32'h13020000;
          16'h01a3 : blkif.rom_rdata <= 32'h9300d000;
          16'h01a4 : blkif.rom_rdata <= 32'h9381b000;
          16'h01a5 : blkif.rom_rdata <= 32'h13830100;
          16'h01a6 : blkif.rom_rdata <= 32'h13021200;
          16'h01a7 : blkif.rom_rdata <= 32'h93022000;
          16'h01a8 : blkif.rom_rdata <= 32'he31652fe;
          16'h01a9 : blkif.rom_rdata <= 32'h930e8001;
          16'h01aa : blkif.rom_rdata <= 32'h130e7003;
          16'h01ab : blkif.rom_rdata <= 32'h6304d301;
          16'h01ac : blkif.rom_rdata <= 32'h6f50c00b;
          16'h01ad : blkif.rom_rdata <= 32'hb7000080;
          16'h01ae : blkif.rom_rdata <= 32'h93804000;
          16'h01af : blkif.rom_rdata <= 32'h13019003;
          16'h01b0 : blkif.rom_rdata <= 32'h23a02000;
          16'h01b1 : blkif.rom_rdata <= 32'h13020000;
          16'h01b2 : blkif.rom_rdata <= 32'h9300d000;
          16'h01b3 : blkif.rom_rdata <= 32'h93819000;
          16'h01b4 : blkif.rom_rdata <= 32'h13000000;
          16'h01b5 : blkif.rom_rdata <= 32'h13000000;
          16'h01b6 : blkif.rom_rdata <= 32'h13830100;
          16'h01b7 : blkif.rom_rdata <= 32'h13021200;
          16'h01b8 : blkif.rom_rdata <= 32'h93022000;
          16'h01b9 : blkif.rom_rdata <= 32'he31252fe;
          16'h01ba : blkif.rom_rdata <= 32'h930e6001;
          16'h01bb : blkif.rom_rdata <= 32'h130e9003;
          16'h01bc : blkif.rom_rdata <= 32'h6304d301;
          16'h01bd : blkif.rom_rdata <= 32'h6f508007;
          16'h01be : blkif.rom_rdata <= 32'hb7000080;
          16'h01bf : blkif.rom_rdata <= 32'h93804000;
          16'h01c0 : blkif.rom_rdata <= 32'h1301a003;
          16'h01c1 : blkif.rom_rdata <= 32'h23a02000;
          16'h01c2 : blkif.rom_rdata <= 32'h13020000;
          16'h01c3 : blkif.rom_rdata <= 32'h9300d000;
          16'h01c4 : blkif.rom_rdata <= 32'h9381b000;
          16'h01c5 : blkif.rom_rdata <= 32'h13021200;
          16'h01c6 : blkif.rom_rdata <= 32'h93022000;
          16'h01c7 : blkif.rom_rdata <= 32'he31852fe;
          16'h01c8 : blkif.rom_rdata <= 32'h930e8001;
          16'h01c9 : blkif.rom_rdata <= 32'h130ea003;
          16'h01ca : blkif.rom_rdata <= 32'h6384d101;
          16'h01cb : blkif.rom_rdata <= 32'h6f500004;
          16'h01cc : blkif.rom_rdata <= 32'hb7000080;
          16'h01cd : blkif.rom_rdata <= 32'h93804000;
          16'h01ce : blkif.rom_rdata <= 32'h1301d003;
          16'h01cf : blkif.rom_rdata <= 32'h23a02000;
          16'h01d0 : blkif.rom_rdata <= 32'h93000002;
          16'h01d1 : blkif.rom_rdata <= 32'h930e0002;
          16'h01d2 : blkif.rom_rdata <= 32'h130ed003;
          16'h01d3 : blkif.rom_rdata <= 32'h6384d001;
          16'h01d4 : blkif.rom_rdata <= 32'h6f50c001;
          16'h01d5 : blkif.rom_rdata <= 32'hb7000080;
          16'h01d6 : blkif.rom_rdata <= 32'h93804000;
          16'h01d7 : blkif.rom_rdata <= 32'h1301e003;
          16'h01d8 : blkif.rom_rdata <= 32'h23a02000;
          16'h01d9 : blkif.rom_rdata <= 32'h93001002;
          16'h01da : blkif.rom_rdata <= 32'h13802003;
          16'h01db : blkif.rom_rdata <= 32'h930e0000;
          16'h01dc : blkif.rom_rdata <= 32'h130ee003;
          16'h01dd : blkif.rom_rdata <= 32'h6304d001;
          16'h01de : blkif.rom_rdata <= 32'h6f40507f;
          16'h01df : blkif.rom_rdata <= 32'hb7000080;
          16'h01e0 : blkif.rom_rdata <= 32'h93804000;
          16'h01e1 : blkif.rom_rdata <= 32'h1301f003;
          16'h01e2 : blkif.rom_rdata <= 32'h23a02000;
          16'h01e3 : blkif.rom_rdata <= 32'hb70001ff;
          16'h01e4 : blkif.rom_rdata <= 32'h938000f0;
          16'h01e5 : blkif.rom_rdata <= 32'h37110f0f;
          16'h01e6 : blkif.rom_rdata <= 32'h1301f1f0;
          16'h01e7 : blkif.rom_rdata <= 32'hb3f12000;
          16'h01e8 : blkif.rom_rdata <= 32'hb71e000f;
          16'h01e9 : blkif.rom_rdata <= 32'h938e0ef0;
          16'h01ea : blkif.rom_rdata <= 32'h130ef003;
          16'h01eb : blkif.rom_rdata <= 32'h6384d101;
          16'h01ec : blkif.rom_rdata <= 32'h6f40d07b;
          16'h01ed : blkif.rom_rdata <= 32'hb7000080;
          16'h01ee : blkif.rom_rdata <= 32'h93804000;
          16'h01ef : blkif.rom_rdata <= 32'h13012004;
          16'h01f0 : blkif.rom_rdata <= 32'h23a02000;
          16'h01f1 : blkif.rom_rdata <= 32'hb7f00ff0;
          16'h01f2 : blkif.rom_rdata <= 32'h9380f000;
          16'h01f3 : blkif.rom_rdata <= 32'h37f1f0f0;
          16'h01f4 : blkif.rom_rdata <= 32'h1301010f;
          16'h01f5 : blkif.rom_rdata <= 32'hb3f12000;
          16'h01f6 : blkif.rom_rdata <= 32'hb7fe00f0;
          16'h01f7 : blkif.rom_rdata <= 32'h130e2004;
          16'h01f8 : blkif.rom_rdata <= 32'h6384d101;
          16'h01f9 : blkif.rom_rdata <= 32'h6f409078;
          16'h01fa : blkif.rom_rdata <= 32'hb7000080;
          16'h01fb : blkif.rom_rdata <= 32'h93804000;
          16'h01fc : blkif.rom_rdata <= 32'h13013004;
          16'h01fd : blkif.rom_rdata <= 32'h23a02000;
          16'h01fe : blkif.rom_rdata <= 32'hb70001ff;
          16'h01ff : blkif.rom_rdata <= 32'h938000f0;
          16'h0200 : blkif.rom_rdata <= 32'h37110f0f;
          16'h0201 : blkif.rom_rdata <= 32'h1301f1f0;
          16'h0202 : blkif.rom_rdata <= 32'hb3f02000;
          16'h0203 : blkif.rom_rdata <= 32'hb71e000f;
          16'h0204 : blkif.rom_rdata <= 32'h938e0ef0;
          16'h0205 : blkif.rom_rdata <= 32'h130e3004;
          16'h0206 : blkif.rom_rdata <= 32'h6384d001;
          16'h0207 : blkif.rom_rdata <= 32'h6f401075;
          16'h0208 : blkif.rom_rdata <= 32'hb7000080;
          16'h0209 : blkif.rom_rdata <= 32'h93804000;
          16'h020a : blkif.rom_rdata <= 32'h13015004;
          16'h020b : blkif.rom_rdata <= 32'h23a02000;
          16'h020c : blkif.rom_rdata <= 32'hb70001ff;
          16'h020d : blkif.rom_rdata <= 32'h938000f0;
          16'h020e : blkif.rom_rdata <= 32'hb3f01000;
          16'h020f : blkif.rom_rdata <= 32'hb70e01ff;
          16'h0210 : blkif.rom_rdata <= 32'h938e0ef0;
          16'h0211 : blkif.rom_rdata <= 32'h130e5004;
          16'h0212 : blkif.rom_rdata <= 32'h6384d001;
          16'h0213 : blkif.rom_rdata <= 32'h6f401072;
          16'h0214 : blkif.rom_rdata <= 32'hb7000080;
          16'h0215 : blkif.rom_rdata <= 32'h93804000;
          16'h0216 : blkif.rom_rdata <= 32'h13016004;
          16'h0217 : blkif.rom_rdata <= 32'h23a02000;
          16'h0218 : blkif.rom_rdata <= 32'h13020000;
          16'h0219 : blkif.rom_rdata <= 32'hb70001ff;
          16'h021a : blkif.rom_rdata <= 32'h938000f0;
          16'h021b : blkif.rom_rdata <= 32'h37110f0f;
          16'h021c : blkif.rom_rdata <= 32'h1301f1f0;
          16'h021d : blkif.rom_rdata <= 32'hb3f12000;
          16'h021e : blkif.rom_rdata <= 32'h13830100;
          16'h021f : blkif.rom_rdata <= 32'h13021200;
          16'h0220 : blkif.rom_rdata <= 32'h93022000;
          16'h0221 : blkif.rom_rdata <= 32'he31052fe;
          16'h0222 : blkif.rom_rdata <= 32'hb71e000f;
          16'h0223 : blkif.rom_rdata <= 32'h938e0ef0;
          16'h0224 : blkif.rom_rdata <= 32'h130e6004;
          16'h0225 : blkif.rom_rdata <= 32'h6304d301;
          16'h0226 : blkif.rom_rdata <= 32'h6f40506d;
          16'h0227 : blkif.rom_rdata <= 32'hb7000080;
          16'h0228 : blkif.rom_rdata <= 32'h93804000;
          16'h0229 : blkif.rom_rdata <= 32'h13018004;
          16'h022a : blkif.rom_rdata <= 32'h23a02000;
          16'h022b : blkif.rom_rdata <= 32'h13020000;
          16'h022c : blkif.rom_rdata <= 32'hb700ff00;
          16'h022d : blkif.rom_rdata <= 32'h9380f00f;
          16'h022e : blkif.rom_rdata <= 32'h37110f0f;
          16'h022f : blkif.rom_rdata <= 32'h1301f1f0;
          16'h0230 : blkif.rom_rdata <= 32'hb3f12000;
          16'h0231 : blkif.rom_rdata <= 32'h13000000;
          16'h0232 : blkif.rom_rdata <= 32'h13000000;
          16'h0233 : blkif.rom_rdata <= 32'h13830100;
          16'h0234 : blkif.rom_rdata <= 32'h13021200;
          16'h0235 : blkif.rom_rdata <= 32'h93022000;
          16'h0236 : blkif.rom_rdata <= 32'he31c52fc;
          16'h0237 : blkif.rom_rdata <= 32'hb70e0f00;
          16'h0238 : blkif.rom_rdata <= 32'h938efe00;
          16'h0239 : blkif.rom_rdata <= 32'h130e8004;
          16'h023a : blkif.rom_rdata <= 32'h6304d301;
          16'h023b : blkif.rom_rdata <= 32'h6f401068;
          16'h023c : blkif.rom_rdata <= 32'hb7000080;
          16'h023d : blkif.rom_rdata <= 32'h93804000;
          16'h023e : blkif.rom_rdata <= 32'h1301f004;
          16'h023f : blkif.rom_rdata <= 32'h23a02000;
          16'h0240 : blkif.rom_rdata <= 32'h13020000;
          16'h0241 : blkif.rom_rdata <= 32'h37110f0f;
          16'h0242 : blkif.rom_rdata <= 32'h1301f1f0;
          16'h0243 : blkif.rom_rdata <= 32'hb70001ff;
          16'h0244 : blkif.rom_rdata <= 32'h938000f0;
          16'h0245 : blkif.rom_rdata <= 32'hb3f12000;
          16'h0246 : blkif.rom_rdata <= 32'h13021200;
          16'h0247 : blkif.rom_rdata <= 32'h93022000;
          16'h0248 : blkif.rom_rdata <= 32'he31252fe;
          16'h0249 : blkif.rom_rdata <= 32'hb71e000f;
          16'h024a : blkif.rom_rdata <= 32'h938e0ef0;
          16'h024b : blkif.rom_rdata <= 32'h130ef004;
          16'h024c : blkif.rom_rdata <= 32'h6384d101;
          16'h024d : blkif.rom_rdata <= 32'h6f409063;
          16'h024e : blkif.rom_rdata <= 32'hb7000080;
          16'h024f : blkif.rom_rdata <= 32'h93804000;
          16'h0250 : blkif.rom_rdata <= 32'h13014005;
          16'h0251 : blkif.rom_rdata <= 32'h23a02000;
          16'h0252 : blkif.rom_rdata <= 32'h13020000;
          16'h0253 : blkif.rom_rdata <= 32'h37110f0f;
          16'h0254 : blkif.rom_rdata <= 32'h1301f1f0;
          16'h0255 : blkif.rom_rdata <= 32'h13000000;
          16'h0256 : blkif.rom_rdata <= 32'h13000000;
          16'h0257 : blkif.rom_rdata <= 32'hb700ff00;
          16'h0258 : blkif.rom_rdata <= 32'h9380f00f;
          16'h0259 : blkif.rom_rdata <= 32'hb3f12000;
          16'h025a : blkif.rom_rdata <= 32'h13021200;
          16'h025b : blkif.rom_rdata <= 32'h93022000;
          16'h025c : blkif.rom_rdata <= 32'he31e52fc;
          16'h025d : blkif.rom_rdata <= 32'hb70e0f00;
          16'h025e : blkif.rom_rdata <= 32'h938efe00;
          16'h025f : blkif.rom_rdata <= 32'h130e4005;
          16'h0260 : blkif.rom_rdata <= 32'h6384d101;
          16'h0261 : blkif.rom_rdata <= 32'h6f40905e;
          16'h0262 : blkif.rom_rdata <= 32'hb7000080;
          16'h0263 : blkif.rom_rdata <= 32'h93804000;
          16'h0264 : blkif.rom_rdata <= 32'h13015005;
          16'h0265 : blkif.rom_rdata <= 32'h23a02000;
          16'h0266 : blkif.rom_rdata <= 32'hb70001ff;
          16'h0267 : blkif.rom_rdata <= 32'h938000f0;
          16'h0268 : blkif.rom_rdata <= 32'h33711000;
          16'h0269 : blkif.rom_rdata <= 32'h930e0000;
          16'h026a : blkif.rom_rdata <= 32'h130e5005;
          16'h026b : blkif.rom_rdata <= 32'h6304d101;
          16'h026c : blkif.rom_rdata <= 32'h6f40d05b;
          16'h026d : blkif.rom_rdata <= 32'hb7000080;
          16'h026e : blkif.rom_rdata <= 32'h93804000;
          16'h026f : blkif.rom_rdata <= 32'h13016005;
          16'h0270 : blkif.rom_rdata <= 32'h23a02000;
          16'h0271 : blkif.rom_rdata <= 32'hb700ff00;
          16'h0272 : blkif.rom_rdata <= 32'h9380f00f;
          16'h0273 : blkif.rom_rdata <= 32'h33f10000;
          16'h0274 : blkif.rom_rdata <= 32'h930e0000;
          16'h0275 : blkif.rom_rdata <= 32'h130e6005;
          16'h0276 : blkif.rom_rdata <= 32'h6304d101;
          16'h0277 : blkif.rom_rdata <= 32'h6f401059;
          16'h0278 : blkif.rom_rdata <= 32'hb7000080;
          16'h0279 : blkif.rom_rdata <= 32'h93804000;
          16'h027a : blkif.rom_rdata <= 32'h13017005;
          16'h027b : blkif.rom_rdata <= 32'h23a02000;
          16'h027c : blkif.rom_rdata <= 32'hb3700000;
          16'h027d : blkif.rom_rdata <= 32'h930e0000;
          16'h027e : blkif.rom_rdata <= 32'h130e7005;
          16'h027f : blkif.rom_rdata <= 32'h6384d001;
          16'h0280 : blkif.rom_rdata <= 32'h6f40d056;
          16'h0281 : blkif.rom_rdata <= 32'hb7000080;
          16'h0282 : blkif.rom_rdata <= 32'h93804000;
          16'h0283 : blkif.rom_rdata <= 32'h13018005;
          16'h0284 : blkif.rom_rdata <= 32'h23a02000;
          16'h0285 : blkif.rom_rdata <= 32'hb7101111;
          16'h0286 : blkif.rom_rdata <= 32'h93801011;
          16'h0287 : blkif.rom_rdata <= 32'h37212222;
          16'h0288 : blkif.rom_rdata <= 32'h13012122;
          16'h0289 : blkif.rom_rdata <= 32'h33f02000;
          16'h028a : blkif.rom_rdata <= 32'h930e0000;
          16'h028b : blkif.rom_rdata <= 32'h130e8005;
          16'h028c : blkif.rom_rdata <= 32'h6304d001;
          16'h028d : blkif.rom_rdata <= 32'h6f409053;
          16'h028e : blkif.rom_rdata <= 32'hb7000080;
          16'h028f : blkif.rom_rdata <= 32'h93804000;
          16'h0290 : blkif.rom_rdata <= 32'h13019005;
          16'h0291 : blkif.rom_rdata <= 32'h23a02000;
          16'h0292 : blkif.rom_rdata <= 32'hb70001ff;
          16'h0293 : blkif.rom_rdata <= 32'h938000f0;
          16'h0294 : blkif.rom_rdata <= 32'h93f1f0f0;
          16'h0295 : blkif.rom_rdata <= 32'hb70e01ff;
          16'h0296 : blkif.rom_rdata <= 32'h938e0ef0;
          16'h0297 : blkif.rom_rdata <= 32'h130e9005;
          16'h0298 : blkif.rom_rdata <= 32'h6384d101;
          16'h0299 : blkif.rom_rdata <= 32'h6f409050;
          16'h029a : blkif.rom_rdata <= 32'hb7000080;
          16'h029b : blkif.rom_rdata <= 32'h93804000;
          16'h029c : blkif.rom_rdata <= 32'h1301b005;
          16'h029d : blkif.rom_rdata <= 32'h23a02000;
          16'h029e : blkif.rom_rdata <= 32'hb700ff00;
          16'h029f : blkif.rom_rdata <= 32'h9380f00f;
          16'h02a0 : blkif.rom_rdata <= 32'h93f1f070;
          16'h02a1 : blkif.rom_rdata <= 32'h930ef000;
          16'h02a2 : blkif.rom_rdata <= 32'h130eb005;
          16'h02a3 : blkif.rom_rdata <= 32'h6384d101;
          16'h02a4 : blkif.rom_rdata <= 32'h6f40d04d;
          16'h02a5 : blkif.rom_rdata <= 32'hb7000080;
          16'h02a6 : blkif.rom_rdata <= 32'h93804000;
          16'h02a7 : blkif.rom_rdata <= 32'h1301c005;
          16'h02a8 : blkif.rom_rdata <= 32'h23a02000;
          16'h02a9 : blkif.rom_rdata <= 32'hb7f00ff0;
          16'h02aa : blkif.rom_rdata <= 32'h9380f000;
          16'h02ab : blkif.rom_rdata <= 32'h93f1000f;
          16'h02ac : blkif.rom_rdata <= 32'h930e0000;
          16'h02ad : blkif.rom_rdata <= 32'h130ec005;
          16'h02ae : blkif.rom_rdata <= 32'h6384d101;
          16'h02af : blkif.rom_rdata <= 32'h6f40104b;
          16'h02b0 : blkif.rom_rdata <= 32'hb7000080;
          16'h02b1 : blkif.rom_rdata <= 32'h93804000;
          16'h02b2 : blkif.rom_rdata <= 32'h1301d005;
          16'h02b3 : blkif.rom_rdata <= 32'h23a02000;
          16'h02b4 : blkif.rom_rdata <= 32'hb70001ff;
          16'h02b5 : blkif.rom_rdata <= 32'h938000f0;
          16'h02b6 : blkif.rom_rdata <= 32'h93f0000f;
          16'h02b7 : blkif.rom_rdata <= 32'h930e0000;
          16'h02b8 : blkif.rom_rdata <= 32'h130ed005;
          16'h02b9 : blkif.rom_rdata <= 32'h6384d001;
          16'h02ba : blkif.rom_rdata <= 32'h6f405048;
          16'h02bb : blkif.rom_rdata <= 32'hb7000080;
          16'h02bc : blkif.rom_rdata <= 32'h93804000;
          16'h02bd : blkif.rom_rdata <= 32'h1301e005;
          16'h02be : blkif.rom_rdata <= 32'h23a02000;
          16'h02bf : blkif.rom_rdata <= 32'h13020000;
          16'h02c0 : blkif.rom_rdata <= 32'hb710f00f;
          16'h02c1 : blkif.rom_rdata <= 32'h938000ff;
          16'h02c2 : blkif.rom_rdata <= 32'h93f1f070;
          16'h02c3 : blkif.rom_rdata <= 32'h13830100;
          16'h02c4 : blkif.rom_rdata <= 32'h13021200;
          16'h02c5 : blkif.rom_rdata <= 32'h93022000;
          16'h02c6 : blkif.rom_rdata <= 32'he31452fe;
          16'h02c7 : blkif.rom_rdata <= 32'h930e0070;
          16'h02c8 : blkif.rom_rdata <= 32'h130ee005;
          16'h02c9 : blkif.rom_rdata <= 32'h6304d301;
          16'h02ca : blkif.rom_rdata <= 32'h6f405044;
          16'h02cb : blkif.rom_rdata <= 32'hb7000080;
          16'h02cc : blkif.rom_rdata <= 32'h93804000;
          16'h02cd : blkif.rom_rdata <= 32'h13010006;
          16'h02ce : blkif.rom_rdata <= 32'h23a02000;
          16'h02cf : blkif.rom_rdata <= 32'h13020000;
          16'h02d0 : blkif.rom_rdata <= 32'hb7f00ff0;
          16'h02d1 : blkif.rom_rdata <= 32'h9380f000;
          16'h02d2 : blkif.rom_rdata <= 32'h93f1f0f0;
          16'h02d3 : blkif.rom_rdata <= 32'h13000000;
          16'h02d4 : blkif.rom_rdata <= 32'h13000000;
          16'h02d5 : blkif.rom_rdata <= 32'h13830100;
          16'h02d6 : blkif.rom_rdata <= 32'h13021200;
          16'h02d7 : blkif.rom_rdata <= 32'h93022000;
          16'h02d8 : blkif.rom_rdata <= 32'he31052fe;
          16'h02d9 : blkif.rom_rdata <= 32'hb7fe0ff0;
          16'h02da : blkif.rom_rdata <= 32'h938efe00;
          16'h02db : blkif.rom_rdata <= 32'h130e0006;
          16'h02dc : blkif.rom_rdata <= 32'h6304d301;
          16'h02dd : blkif.rom_rdata <= 32'h6f40903f;
          16'h02de : blkif.rom_rdata <= 32'hb7000080;
          16'h02df : blkif.rom_rdata <= 32'h93804000;
          16'h02e0 : blkif.rom_rdata <= 32'h13014006;
          16'h02e1 : blkif.rom_rdata <= 32'h23a02000;
          16'h02e2 : blkif.rom_rdata <= 32'h9370000f;
          16'h02e3 : blkif.rom_rdata <= 32'h930e0000;
          16'h02e4 : blkif.rom_rdata <= 32'h130e4006;
          16'h02e5 : blkif.rom_rdata <= 32'h6384d001;
          16'h02e6 : blkif.rom_rdata <= 32'h6f40503d;
          16'h02e7 : blkif.rom_rdata <= 32'hb7000080;
          16'h02e8 : blkif.rom_rdata <= 32'h93804000;
          16'h02e9 : blkif.rom_rdata <= 32'h13015006;
          16'h02ea : blkif.rom_rdata <= 32'h23a02000;
          16'h02eb : blkif.rom_rdata <= 32'hb700ff00;
          16'h02ec : blkif.rom_rdata <= 32'h9380f00f;
          16'h02ed : blkif.rom_rdata <= 32'h13f0f070;
          16'h02ee : blkif.rom_rdata <= 32'h930e0000;
          16'h02ef : blkif.rom_rdata <= 32'h130e5006;
          16'h02f0 : blkif.rom_rdata <= 32'h6304d001;
          16'h02f1 : blkif.rom_rdata <= 32'h6f40903a;
          16'h02f2 : blkif.rom_rdata <= 32'hb7000080;
          16'h02f3 : blkif.rom_rdata <= 32'h93804000;
          16'h02f4 : blkif.rom_rdata <= 32'h13016006;
          16'h02f5 : blkif.rom_rdata <= 32'h23a02000;
          16'h02f6 : blkif.rom_rdata <= 32'h17250000;
          16'h02f7 : blkif.rom_rdata <= 32'h1305c571;
          16'h02f8 : blkif.rom_rdata <= 32'hef054000;
          16'h02f9 : blkif.rom_rdata <= 32'h3305b540;
          16'h02fa : blkif.rom_rdata <= 32'hb72e0000;
          16'h02fb : blkif.rom_rdata <= 32'h938e0e71;
          16'h02fc : blkif.rom_rdata <= 32'h130e6006;
          16'h02fd : blkif.rom_rdata <= 32'h6304d501;
          16'h02fe : blkif.rom_rdata <= 32'h6f405037;
          16'h02ff : blkif.rom_rdata <= 32'hb7000080;
          16'h0300 : blkif.rom_rdata <= 32'h93804000;
          16'h0301 : blkif.rom_rdata <= 32'h13017006;
          16'h0302 : blkif.rom_rdata <= 32'h23a02000;
          16'h0303 : blkif.rom_rdata <= 32'h13000000;
          16'h0304 : blkif.rom_rdata <= 32'h17e5ffff;
          16'h0305 : blkif.rom_rdata <= 32'h1305c58f;
          16'h0306 : blkif.rom_rdata <= 32'hef054000;
          16'h0307 : blkif.rom_rdata <= 32'h3305b540;
          16'h0308 : blkif.rom_rdata <= 32'hb7eeffff;
          16'h0309 : blkif.rom_rdata <= 32'h938e0e8f;
          16'h030a : blkif.rom_rdata <= 32'h130e7006;
          16'h030b : blkif.rom_rdata <= 32'h6304d501;
          16'h030c : blkif.rom_rdata <= 32'h6f40d033;
          16'h030d : blkif.rom_rdata <= 32'h130e8006;
          16'h030e : blkif.rom_rdata <= 32'h93000000;
          16'h030f : blkif.rom_rdata <= 32'h13010000;
          16'h0310 : blkif.rom_rdata <= 32'h63882000;
          16'h0311 : blkif.rom_rdata <= 32'h6304c001;
          16'h0312 : blkif.rom_rdata <= 32'h6f405032;
          16'h0313 : blkif.rom_rdata <= 32'h6318c001;
          16'h0314 : blkif.rom_rdata <= 32'he38e20fe;
          16'h0315 : blkif.rom_rdata <= 32'h6304c001;
          16'h0316 : blkif.rom_rdata <= 32'h6f405031;
          16'h0317 : blkif.rom_rdata <= 32'h130ea006;
          16'h0318 : blkif.rom_rdata <= 32'h9300f0ff;
          16'h0319 : blkif.rom_rdata <= 32'h1301f0ff;
          16'h031a : blkif.rom_rdata <= 32'h63882000;
          16'h031b : blkif.rom_rdata <= 32'h6304c001;
          16'h031c : blkif.rom_rdata <= 32'h6f40d02f;
          16'h031d : blkif.rom_rdata <= 32'h6318c001;
          16'h031e : blkif.rom_rdata <= 32'he38e20fe;
          16'h031f : blkif.rom_rdata <= 32'h6304c001;
          16'h0320 : blkif.rom_rdata <= 32'h6f40d02e;
          16'h0321 : blkif.rom_rdata <= 32'h130ef006;
          16'h0322 : blkif.rom_rdata <= 32'h13020000;
          16'h0323 : blkif.rom_rdata <= 32'h93000000;
          16'h0324 : blkif.rom_rdata <= 32'h1301f0ff;
          16'h0325 : blkif.rom_rdata <= 32'h63942000;
          16'h0326 : blkif.rom_rdata <= 32'h6f40502d;
          16'h0327 : blkif.rom_rdata <= 32'h13021200;
          16'h0328 : blkif.rom_rdata <= 32'h93022000;
          16'h0329 : blkif.rom_rdata <= 32'he31452fe;
          16'h032a : blkif.rom_rdata <= 32'h130e4007;
          16'h032b : blkif.rom_rdata <= 32'h13020000;
          16'h032c : blkif.rom_rdata <= 32'h93000000;
          16'h032d : blkif.rom_rdata <= 32'h13000000;
          16'h032e : blkif.rom_rdata <= 32'h13000000;
          16'h032f : blkif.rom_rdata <= 32'h1301f0ff;
          16'h0330 : blkif.rom_rdata <= 32'h63942000;
          16'h0331 : blkif.rom_rdata <= 32'h6f40902a;
          16'h0332 : blkif.rom_rdata <= 32'h13021200;
          16'h0333 : blkif.rom_rdata <= 32'h93022000;
          16'h0334 : blkif.rom_rdata <= 32'he31052fe;
          16'h0335 : blkif.rom_rdata <= 32'h130e5007;
          16'h0336 : blkif.rom_rdata <= 32'h13020000;
          16'h0337 : blkif.rom_rdata <= 32'h93000000;
          16'h0338 : blkif.rom_rdata <= 32'h1301f0ff;
          16'h0339 : blkif.rom_rdata <= 32'h63942000;
          16'h033a : blkif.rom_rdata <= 32'h6f405028;
          16'h033b : blkif.rom_rdata <= 32'h13021200;
          16'h033c : blkif.rom_rdata <= 32'h93022000;
          16'h033d : blkif.rom_rdata <= 32'he31452fe;
          16'h033e : blkif.rom_rdata <= 32'h130ea007;
          16'h033f : blkif.rom_rdata <= 32'h13020000;
          16'h0340 : blkif.rom_rdata <= 32'h93000000;
          16'h0341 : blkif.rom_rdata <= 32'h13000000;
          16'h0342 : blkif.rom_rdata <= 32'h13000000;
          16'h0343 : blkif.rom_rdata <= 32'h1301f0ff;
          16'h0344 : blkif.rom_rdata <= 32'h63942000;
          16'h0345 : blkif.rom_rdata <= 32'h6f409025;
          16'h0346 : blkif.rom_rdata <= 32'h13021200;
          16'h0347 : blkif.rom_rdata <= 32'h93022000;
          16'h0348 : blkif.rom_rdata <= 32'he31052fe;
          16'h0349 : blkif.rom_rdata <= 32'hb7000080;
          16'h034a : blkif.rom_rdata <= 32'h93804000;
          16'h034b : blkif.rom_rdata <= 32'h1301b007;
          16'h034c : blkif.rom_rdata <= 32'h23a02000;
          16'h034d : blkif.rom_rdata <= 32'h93001000;
          16'h034e : blkif.rom_rdata <= 32'h630a0000;
          16'h034f : blkif.rom_rdata <= 32'h93801000;
          16'h0350 : blkif.rom_rdata <= 32'h93801000;
          16'h0351 : blkif.rom_rdata <= 32'h93801000;
          16'h0352 : blkif.rom_rdata <= 32'h93801000;
          16'h0353 : blkif.rom_rdata <= 32'h93801000;
          16'h0354 : blkif.rom_rdata <= 32'h93801000;
          16'h0355 : blkif.rom_rdata <= 32'h930e3000;
          16'h0356 : blkif.rom_rdata <= 32'h130eb007;
          16'h0357 : blkif.rom_rdata <= 32'h6384d001;
          16'h0358 : blkif.rom_rdata <= 32'h6f40d020;
          16'h0359 : blkif.rom_rdata <= 32'h130ec007;
          16'h035a : blkif.rom_rdata <= 32'h93000000;
          16'h035b : blkif.rom_rdata <= 32'h13010000;
          16'h035c : blkif.rom_rdata <= 32'h63d82000;
          16'h035d : blkif.rom_rdata <= 32'h6304c001;
          16'h035e : blkif.rom_rdata <= 32'h6f40501f;
          16'h035f : blkif.rom_rdata <= 32'h6318c001;
          16'h0360 : blkif.rom_rdata <= 32'he3de20fe;
          16'h0361 : blkif.rom_rdata <= 32'h6304c001;
          16'h0362 : blkif.rom_rdata <= 32'h6f40501e;
          16'h0363 : blkif.rom_rdata <= 32'h130e1008;
          16'h0364 : blkif.rom_rdata <= 32'h9300f0ff;
          16'h0365 : blkif.rom_rdata <= 32'h1301e0ff;
          16'h0366 : blkif.rom_rdata <= 32'h63d82000;
          16'h0367 : blkif.rom_rdata <= 32'h6304c001;
          16'h0368 : blkif.rom_rdata <= 32'h6f40d01c;
          16'h0369 : blkif.rom_rdata <= 32'h6318c001;
          16'h036a : blkif.rom_rdata <= 32'he3de20fe;
          16'h036b : blkif.rom_rdata <= 32'h6304c001;
          16'h036c : blkif.rom_rdata <= 32'h6f40d01b;
          16'h036d : blkif.rom_rdata <= 32'h130e2008;
          16'h036e : blkif.rom_rdata <= 32'h93000000;
          16'h036f : blkif.rom_rdata <= 32'h13011000;
          16'h0370 : blkif.rom_rdata <= 32'h63d42000;
          16'h0371 : blkif.rom_rdata <= 32'h6316c001;
          16'h0372 : blkif.rom_rdata <= 32'h6304c001;
          16'h0373 : blkif.rom_rdata <= 32'h6f40101a;
          16'h0374 : blkif.rom_rdata <= 32'he3dc20fe;
          16'h0375 : blkif.rom_rdata <= 32'h130e5008;
          16'h0376 : blkif.rom_rdata <= 32'h9300e0ff;
          16'h0377 : blkif.rom_rdata <= 32'h13011000;
          16'h0378 : blkif.rom_rdata <= 32'h63d42000;
          16'h0379 : blkif.rom_rdata <= 32'h6316c001;
          16'h037a : blkif.rom_rdata <= 32'h6304c001;
          16'h037b : blkif.rom_rdata <= 32'h6f401018;
          16'h037c : blkif.rom_rdata <= 32'he3dc20fe;
          16'h037d : blkif.rom_rdata <= 32'h130eb008;
          16'h037e : blkif.rom_rdata <= 32'h13020000;
          16'h037f : blkif.rom_rdata <= 32'h9300f0ff;
          16'h0380 : blkif.rom_rdata <= 32'h13000000;
          16'h0381 : blkif.rom_rdata <= 32'h13000000;
          16'h0382 : blkif.rom_rdata <= 32'h13010000;
          16'h0383 : blkif.rom_rdata <= 32'h63c42000;
          16'h0384 : blkif.rom_rdata <= 32'h6f40d015;
          16'h0385 : blkif.rom_rdata <= 32'h13021200;
          16'h0386 : blkif.rom_rdata <= 32'h93022000;
          16'h0387 : blkif.rom_rdata <= 32'he31052fe;
          16'h0388 : blkif.rom_rdata <= 32'h130ec008;
          16'h0389 : blkif.rom_rdata <= 32'h13020000;
          16'h038a : blkif.rom_rdata <= 32'h9300f0ff;
          16'h038b : blkif.rom_rdata <= 32'h13010000;
          16'h038c : blkif.rom_rdata <= 32'h63c42000;
          16'h038d : blkif.rom_rdata <= 32'h6f409013;
          16'h038e : blkif.rom_rdata <= 32'h13021200;
          16'h038f : blkif.rom_rdata <= 32'h93022000;
          16'h0390 : blkif.rom_rdata <= 32'he31452fe;
          16'h0391 : blkif.rom_rdata <= 32'h130e1009;
          16'h0392 : blkif.rom_rdata <= 32'h13020000;
          16'h0393 : blkif.rom_rdata <= 32'h9300f0ff;
          16'h0394 : blkif.rom_rdata <= 32'h13000000;
          16'h0395 : blkif.rom_rdata <= 32'h13000000;
          16'h0396 : blkif.rom_rdata <= 32'h13010000;
          16'h0397 : blkif.rom_rdata <= 32'h63c42000;
          16'h0398 : blkif.rom_rdata <= 32'h6f40d010;
          16'h0399 : blkif.rom_rdata <= 32'h13021200;
          16'h039a : blkif.rom_rdata <= 32'h93022000;
          16'h039b : blkif.rom_rdata <= 32'he31052fe;
          16'h039c : blkif.rom_rdata <= 32'hb7000080;
          16'h039d : blkif.rom_rdata <= 32'h93804000;
          16'h039e : blkif.rom_rdata <= 32'h13012009;
          16'h039f : blkif.rom_rdata <= 32'h23a02000;
          16'h03a0 : blkif.rom_rdata <= 32'h93001000;
          16'h03a1 : blkif.rom_rdata <= 32'h63da0000;
          16'h03a2 : blkif.rom_rdata <= 32'h93801000;
          16'h03a3 : blkif.rom_rdata <= 32'h93801000;
          16'h03a4 : blkif.rom_rdata <= 32'h93801000;
          16'h03a5 : blkif.rom_rdata <= 32'h93801000;
          16'h03a6 : blkif.rom_rdata <= 32'h93801000;
          16'h03a7 : blkif.rom_rdata <= 32'h93801000;
          16'h03a8 : blkif.rom_rdata <= 32'h930e3000;
          16'h03a9 : blkif.rom_rdata <= 32'h130e2009;
          16'h03aa : blkif.rom_rdata <= 32'h6384d001;
          16'h03ab : blkif.rom_rdata <= 32'h6f40100c;
          16'h03ac : blkif.rom_rdata <= 32'h130e3009;
          16'h03ad : blkif.rom_rdata <= 32'h93000000;
          16'h03ae : blkif.rom_rdata <= 32'h13010000;
          16'h03af : blkif.rom_rdata <= 32'h63f82000;
          16'h03b0 : blkif.rom_rdata <= 32'h6304c001;
          16'h03b1 : blkif.rom_rdata <= 32'h6f40900a;
          16'h03b2 : blkif.rom_rdata <= 32'h6318c001;
          16'h03b3 : blkif.rom_rdata <= 32'he3fe20fe;
          16'h03b4 : blkif.rom_rdata <= 32'h6304c001;
          16'h03b5 : blkif.rom_rdata <= 32'h6f409009;
          16'h03b6 : blkif.rom_rdata <= 32'h130e8009;
          16'h03b7 : blkif.rom_rdata <= 32'h9300f0ff;
          16'h03b8 : blkif.rom_rdata <= 32'h13010000;
          16'h03b9 : blkif.rom_rdata <= 32'h63f82000;
          16'h03ba : blkif.rom_rdata <= 32'h6304c001;
          16'h03bb : blkif.rom_rdata <= 32'h6f401008;
          16'h03bc : blkif.rom_rdata <= 32'h6318c001;
          16'h03bd : blkif.rom_rdata <= 32'he3fe20fe;
          16'h03be : blkif.rom_rdata <= 32'h6304c001;
          16'h03bf : blkif.rom_rdata <= 32'h6f401007;
          16'h03c0 : blkif.rom_rdata <= 32'h130e9009;
          16'h03c1 : blkif.rom_rdata <= 32'h93000000;
          16'h03c2 : blkif.rom_rdata <= 32'h13011000;
          16'h03c3 : blkif.rom_rdata <= 32'h63f42000;
          16'h03c4 : blkif.rom_rdata <= 32'h6316c001;
          16'h03c5 : blkif.rom_rdata <= 32'h6304c001;
          16'h03c6 : blkif.rom_rdata <= 32'h6f405005;
          16'h03c7 : blkif.rom_rdata <= 32'he3fc20fe;
          16'h03c8 : blkif.rom_rdata <= 32'h130ed009;
          16'h03c9 : blkif.rom_rdata <= 32'h13020000;
          16'h03ca : blkif.rom_rdata <= 32'hb70000f0;
          16'h03cb : blkif.rom_rdata <= 32'h9380f0ff;
          16'h03cc : blkif.rom_rdata <= 32'h370100f0;
          16'h03cd : blkif.rom_rdata <= 32'h63e42000;
          16'h03ce : blkif.rom_rdata <= 32'h6f405003;
          16'h03cf : blkif.rom_rdata <= 32'h13021200;
          16'h03d0 : blkif.rom_rdata <= 32'h93022000;
          16'h03d1 : blkif.rom_rdata <= 32'he31252fe;
          16'h03d2 : blkif.rom_rdata <= 32'h130e800a;
          16'h03d3 : blkif.rom_rdata <= 32'h13020000;
          16'h03d4 : blkif.rom_rdata <= 32'hb70000f0;
          16'h03d5 : blkif.rom_rdata <= 32'h9380f0ff;
          16'h03d6 : blkif.rom_rdata <= 32'h13000000;
          16'h03d7 : blkif.rom_rdata <= 32'h13000000;
          16'h03d8 : blkif.rom_rdata <= 32'h370100f0;
          16'h03d9 : blkif.rom_rdata <= 32'h63e42000;
          16'h03da : blkif.rom_rdata <= 32'h6f405000;
          16'h03db : blkif.rom_rdata <= 32'h13021200;
          16'h03dc : blkif.rom_rdata <= 32'h93022000;
          16'h03dd : blkif.rom_rdata <= 32'he31e52fc;
          16'h03de : blkif.rom_rdata <= 32'hb7000080;
          16'h03df : blkif.rom_rdata <= 32'h93804000;
          16'h03e0 : blkif.rom_rdata <= 32'h1301900a;
          16'h03e1 : blkif.rom_rdata <= 32'h23a02000;
          16'h03e2 : blkif.rom_rdata <= 32'h93001000;
          16'h03e3 : blkif.rom_rdata <= 32'h63fa0000;
          16'h03e4 : blkif.rom_rdata <= 32'h93801000;
          16'h03e5 : blkif.rom_rdata <= 32'h93801000;
          16'h03e6 : blkif.rom_rdata <= 32'h93801000;
          16'h03e7 : blkif.rom_rdata <= 32'h93801000;
          16'h03e8 : blkif.rom_rdata <= 32'h93801000;
          16'h03e9 : blkif.rom_rdata <= 32'h93801000;
          16'h03ea : blkif.rom_rdata <= 32'h930e3000;
          16'h03eb : blkif.rom_rdata <= 32'h130e900a;
          16'h03ec : blkif.rom_rdata <= 32'h6384d001;
          16'h03ed : blkif.rom_rdata <= 32'h6f40807b;
          16'h03ee : blkif.rom_rdata <= 32'h130ea00a;
          16'h03ef : blkif.rom_rdata <= 32'h93000000;
          16'h03f0 : blkif.rom_rdata <= 32'h13011000;
          16'h03f1 : blkif.rom_rdata <= 32'h63c82000;
          16'h03f2 : blkif.rom_rdata <= 32'h6304c001;
          16'h03f3 : blkif.rom_rdata <= 32'h6f40007a;
          16'h03f4 : blkif.rom_rdata <= 32'h6318c001;
          16'h03f5 : blkif.rom_rdata <= 32'he3ce20fe;
          16'h03f6 : blkif.rom_rdata <= 32'h6304c001;
          16'h03f7 : blkif.rom_rdata <= 32'h6f400079;
          16'h03f8 : blkif.rom_rdata <= 32'h130ec00a;
          16'h03f9 : blkif.rom_rdata <= 32'h9300e0ff;
          16'h03fa : blkif.rom_rdata <= 32'h1301f0ff;
          16'h03fb : blkif.rom_rdata <= 32'h63c82000;
          16'h03fc : blkif.rom_rdata <= 32'h6304c001;
          16'h03fd : blkif.rom_rdata <= 32'h6f408077;
          16'h03fe : blkif.rom_rdata <= 32'h6318c001;
          16'h03ff : blkif.rom_rdata <= 32'he3ce20fe;
          16'h0400 : blkif.rom_rdata <= 32'h6304c001;
          16'h0401 : blkif.rom_rdata <= 32'h6f408076;
          16'h0402 : blkif.rom_rdata <= 32'h130ed00a;
          16'h0403 : blkif.rom_rdata <= 32'h93001000;
          16'h0404 : blkif.rom_rdata <= 32'h13010000;
          16'h0405 : blkif.rom_rdata <= 32'h63c42000;
          16'h0406 : blkif.rom_rdata <= 32'h6316c001;
          16'h0407 : blkif.rom_rdata <= 32'h6304c001;
          16'h0408 : blkif.rom_rdata <= 32'h6f40c074;
          16'h0409 : blkif.rom_rdata <= 32'he3cc20fe;
          16'h040a : blkif.rom_rdata <= 32'h130e000b;
          16'h040b : blkif.rom_rdata <= 32'h93001000;
          16'h040c : blkif.rom_rdata <= 32'h1301e0ff;
          16'h040d : blkif.rom_rdata <= 32'h63c42000;
          16'h040e : blkif.rom_rdata <= 32'h6316c001;
          16'h040f : blkif.rom_rdata <= 32'h6304c001;
          16'h0410 : blkif.rom_rdata <= 32'h6f40c072;
          16'h0411 : blkif.rom_rdata <= 32'he3cc20fe;
          16'h0412 : blkif.rom_rdata <= 32'h130e100b;
          16'h0413 : blkif.rom_rdata <= 32'h13020000;
          16'h0414 : blkif.rom_rdata <= 32'h93000000;
          16'h0415 : blkif.rom_rdata <= 32'h1301f0ff;
          16'h0416 : blkif.rom_rdata <= 32'h63d42000;
          16'h0417 : blkif.rom_rdata <= 32'h6f400071;
          16'h0418 : blkif.rom_rdata <= 32'h13021200;
          16'h0419 : blkif.rom_rdata <= 32'h93022000;
          16'h041a : blkif.rom_rdata <= 32'he31452fe;
          16'h041b : blkif.rom_rdata <= 32'h130ec00b;
          16'h041c : blkif.rom_rdata <= 32'h13020000;
          16'h041d : blkif.rom_rdata <= 32'h93000000;
          16'h041e : blkif.rom_rdata <= 32'h13000000;
          16'h041f : blkif.rom_rdata <= 32'h13000000;
          16'h0420 : blkif.rom_rdata <= 32'h1301f0ff;
          16'h0421 : blkif.rom_rdata <= 32'h63d42000;
          16'h0422 : blkif.rom_rdata <= 32'h6f40406e;
          16'h0423 : blkif.rom_rdata <= 32'h13021200;
          16'h0424 : blkif.rom_rdata <= 32'h93022000;
          16'h0425 : blkif.rom_rdata <= 32'he31052fe;
          16'h0426 : blkif.rom_rdata <= 32'hb7000080;
          16'h0427 : blkif.rom_rdata <= 32'h93804000;
          16'h0428 : blkif.rom_rdata <= 32'h1301d00b;
          16'h0429 : blkif.rom_rdata <= 32'h23a02000;
          16'h042a : blkif.rom_rdata <= 32'h93001000;
          16'h042b : blkif.rom_rdata <= 32'h634a1000;
          16'h042c : blkif.rom_rdata <= 32'h93801000;
          16'h042d : blkif.rom_rdata <= 32'h93801000;
          16'h042e : blkif.rom_rdata <= 32'h93801000;
          16'h042f : blkif.rom_rdata <= 32'h93801000;
          16'h0430 : blkif.rom_rdata <= 32'h93801000;
          16'h0431 : blkif.rom_rdata <= 32'h93801000;
          16'h0432 : blkif.rom_rdata <= 32'h930e3000;
          16'h0433 : blkif.rom_rdata <= 32'h130ed00b;
          16'h0434 : blkif.rom_rdata <= 32'h6384d001;
          16'h0435 : blkif.rom_rdata <= 32'h6f408069;
          16'h0436 : blkif.rom_rdata <= 32'h130ee00b;
          16'h0437 : blkif.rom_rdata <= 32'h93000000;
          16'h0438 : blkif.rom_rdata <= 32'h13011000;
          16'h0439 : blkif.rom_rdata <= 32'h63e82000;
          16'h043a : blkif.rom_rdata <= 32'h6304c001;
          16'h043b : blkif.rom_rdata <= 32'h6f400068;
          16'h043c : blkif.rom_rdata <= 32'h6318c001;
          16'h043d : blkif.rom_rdata <= 32'he3ee20fe;
          16'h043e : blkif.rom_rdata <= 32'h6304c001;
          16'h043f : blkif.rom_rdata <= 32'h6f400067;
          16'h0440 : blkif.rom_rdata <= 32'h130e000c;
          16'h0441 : blkif.rom_rdata <= 32'h93000000;
          16'h0442 : blkif.rom_rdata <= 32'h1301f0ff;
          16'h0443 : blkif.rom_rdata <= 32'h63e82000;
          16'h0444 : blkif.rom_rdata <= 32'h6304c001;
          16'h0445 : blkif.rom_rdata <= 32'h6f408065;
          16'h0446 : blkif.rom_rdata <= 32'h6318c001;
          16'h0447 : blkif.rom_rdata <= 32'he3ee20fe;
          16'h0448 : blkif.rom_rdata <= 32'h6304c001;
          16'h0449 : blkif.rom_rdata <= 32'h6f408064;
          16'h044a : blkif.rom_rdata <= 32'h130e500c;
          16'h044b : blkif.rom_rdata <= 32'h13020000;
          16'h044c : blkif.rom_rdata <= 32'hb70000f0;
          16'h044d : blkif.rom_rdata <= 32'h370100f0;
          16'h044e : blkif.rom_rdata <= 32'h1301f1ff;
          16'h044f : blkif.rom_rdata <= 32'h63f42000;
          16'h0450 : blkif.rom_rdata <= 32'h6f40c062;
          16'h0451 : blkif.rom_rdata <= 32'h13021200;
          16'h0452 : blkif.rom_rdata <= 32'h93022000;
          16'h0453 : blkif.rom_rdata <= 32'he31252fe;
          16'h0454 : blkif.rom_rdata <= 32'h130ea00c;
          16'h0455 : blkif.rom_rdata <= 32'h13020000;
          16'h0456 : blkif.rom_rdata <= 32'hb70000f0;
          16'h0457 : blkif.rom_rdata <= 32'h13000000;
          16'h0458 : blkif.rom_rdata <= 32'h13000000;
          16'h0459 : blkif.rom_rdata <= 32'h370100f0;
          16'h045a : blkif.rom_rdata <= 32'h1301f1ff;
          16'h045b : blkif.rom_rdata <= 32'h63f42000;
          16'h045c : blkif.rom_rdata <= 32'h6f40c05f;
          16'h045d : blkif.rom_rdata <= 32'h13021200;
          16'h045e : blkif.rom_rdata <= 32'h93022000;
          16'h045f : blkif.rom_rdata <= 32'he31e52fc;
          16'h0460 : blkif.rom_rdata <= 32'h130eb00c;
          16'h0461 : blkif.rom_rdata <= 32'h13020000;
          16'h0462 : blkif.rom_rdata <= 32'hb70000f0;
          16'h0463 : blkif.rom_rdata <= 32'h370100f0;
          16'h0464 : blkif.rom_rdata <= 32'h1301f1ff;
          16'h0465 : blkif.rom_rdata <= 32'h63f42000;
          16'h0466 : blkif.rom_rdata <= 32'h6f40405d;
          16'h0467 : blkif.rom_rdata <= 32'h13021200;
          16'h0468 : blkif.rom_rdata <= 32'h93022000;
          16'h0469 : blkif.rom_rdata <= 32'he31252fe;
          16'h046a : blkif.rom_rdata <= 32'h130e000d;
          16'h046b : blkif.rom_rdata <= 32'h13020000;
          16'h046c : blkif.rom_rdata <= 32'hb70000f0;
          16'h046d : blkif.rom_rdata <= 32'h13000000;
          16'h046e : blkif.rom_rdata <= 32'h13000000;
          16'h046f : blkif.rom_rdata <= 32'h370100f0;
          16'h0470 : blkif.rom_rdata <= 32'h1301f1ff;
          16'h0471 : blkif.rom_rdata <= 32'h63f42000;
          16'h0472 : blkif.rom_rdata <= 32'h6f40405a;
          16'h0473 : blkif.rom_rdata <= 32'h13021200;
          16'h0474 : blkif.rom_rdata <= 32'h93022000;
          16'h0475 : blkif.rom_rdata <= 32'he31e52fc;
          16'h0476 : blkif.rom_rdata <= 32'hb7000080;
          16'h0477 : blkif.rom_rdata <= 32'h93804000;
          16'h0478 : blkif.rom_rdata <= 32'h1301100d;
          16'h0479 : blkif.rom_rdata <= 32'h23a02000;
          16'h047a : blkif.rom_rdata <= 32'h93001000;
          16'h047b : blkif.rom_rdata <= 32'h636a1000;
          16'h047c : blkif.rom_rdata <= 32'h93801000;
          16'h047d : blkif.rom_rdata <= 32'h93801000;
          16'h047e : blkif.rom_rdata <= 32'h93801000;
          16'h047f : blkif.rom_rdata <= 32'h93801000;
          16'h0480 : blkif.rom_rdata <= 32'h93801000;
          16'h0481 : blkif.rom_rdata <= 32'h93801000;
          16'h0482 : blkif.rom_rdata <= 32'h930e3000;
          16'h0483 : blkif.rom_rdata <= 32'h130e100d;
          16'h0484 : blkif.rom_rdata <= 32'h6384d001;
          16'h0485 : blkif.rom_rdata <= 32'h6f408055;
          16'h0486 : blkif.rom_rdata <= 32'h130e200d;
          16'h0487 : blkif.rom_rdata <= 32'h93000000;
          16'h0488 : blkif.rom_rdata <= 32'h13011000;
          16'h0489 : blkif.rom_rdata <= 32'h63982000;
          16'h048a : blkif.rom_rdata <= 32'h6304c001;
          16'h048b : blkif.rom_rdata <= 32'h6f400054;
          16'h048c : blkif.rom_rdata <= 32'h6318c001;
          16'h048d : blkif.rom_rdata <= 32'he39e20fe;
          16'h048e : blkif.rom_rdata <= 32'h6304c001;
          16'h048f : blkif.rom_rdata <= 32'h6f400053;
          16'h0490 : blkif.rom_rdata <= 32'h130e500d;
          16'h0491 : blkif.rom_rdata <= 32'h93001000;
          16'h0492 : blkif.rom_rdata <= 32'h1301f0ff;
          16'h0493 : blkif.rom_rdata <= 32'h63982000;
          16'h0494 : blkif.rom_rdata <= 32'h6304c001;
          16'h0495 : blkif.rom_rdata <= 32'h6f408051;
          16'h0496 : blkif.rom_rdata <= 32'h6318c001;
          16'h0497 : blkif.rom_rdata <= 32'he39e20fe;
          16'h0498 : blkif.rom_rdata <= 32'h6304c001;
          16'h0499 : blkif.rom_rdata <= 32'h6f408050;
          16'h049a : blkif.rom_rdata <= 32'h130e600d;
          16'h049b : blkif.rom_rdata <= 32'h93000000;
          16'h049c : blkif.rom_rdata <= 32'h13010000;
          16'h049d : blkif.rom_rdata <= 32'h63942000;
          16'h049e : blkif.rom_rdata <= 32'h6316c001;
          16'h049f : blkif.rom_rdata <= 32'h6304c001;
          16'h04a0 : blkif.rom_rdata <= 32'h6f40c04e;
          16'h04a1 : blkif.rom_rdata <= 32'he39c20fe;
          16'h04a2 : blkif.rom_rdata <= 32'h130e800d;
          16'h04a3 : blkif.rom_rdata <= 32'h9300f0ff;
          16'h04a4 : blkif.rom_rdata <= 32'h1301f0ff;
          16'h04a5 : blkif.rom_rdata <= 32'h63942000;
          16'h04a6 : blkif.rom_rdata <= 32'h6316c001;
          16'h04a7 : blkif.rom_rdata <= 32'h6304c001;
          16'h04a8 : blkif.rom_rdata <= 32'h6f40c04c;
          16'h04a9 : blkif.rom_rdata <= 32'he39c20fe;
          16'h04aa : blkif.rom_rdata <= 32'h130ef00d;
          16'h04ab : blkif.rom_rdata <= 32'h13020000;
          16'h04ac : blkif.rom_rdata <= 32'h93000000;
          16'h04ad : blkif.rom_rdata <= 32'h13010000;
          16'h04ae : blkif.rom_rdata <= 32'h63842000;
          16'h04af : blkif.rom_rdata <= 32'h6f40004b;
          16'h04b0 : blkif.rom_rdata <= 32'h13021200;
          16'h04b1 : blkif.rom_rdata <= 32'h93022000;
          16'h04b2 : blkif.rom_rdata <= 32'he31452fe;
          16'h04b3 : blkif.rom_rdata <= 32'h130e000e;
          16'h04b4 : blkif.rom_rdata <= 32'h13020000;
          16'h04b5 : blkif.rom_rdata <= 32'h93000000;
          16'h04b6 : blkif.rom_rdata <= 32'h13010000;
          16'h04b7 : blkif.rom_rdata <= 32'h13000000;
          16'h04b8 : blkif.rom_rdata <= 32'h63842000;
          16'h04b9 : blkif.rom_rdata <= 32'h6f408048;
          16'h04ba : blkif.rom_rdata <= 32'h13021200;
          16'h04bb : blkif.rom_rdata <= 32'h93022000;
          16'h04bc : blkif.rom_rdata <= 32'he31252fe;
          16'h04bd : blkif.rom_rdata <= 32'h130e400e;
          16'h04be : blkif.rom_rdata <= 32'h13020000;
          16'h04bf : blkif.rom_rdata <= 32'h93000000;
          16'h04c0 : blkif.rom_rdata <= 32'h13000000;
          16'h04c1 : blkif.rom_rdata <= 32'h13000000;
          16'h04c2 : blkif.rom_rdata <= 32'h13010000;
          16'h04c3 : blkif.rom_rdata <= 32'h63842000;
          16'h04c4 : blkif.rom_rdata <= 32'h6f40c045;
          16'h04c5 : blkif.rom_rdata <= 32'h13021200;
          16'h04c6 : blkif.rom_rdata <= 32'h93022000;
          16'h04c7 : blkif.rom_rdata <= 32'he31052fe;
          16'h04c8 : blkif.rom_rdata <= 32'hb7000080;
          16'h04c9 : blkif.rom_rdata <= 32'h93804000;
          16'h04ca : blkif.rom_rdata <= 32'h1301500e;
          16'h04cb : blkif.rom_rdata <= 32'h23a02000;
          16'h04cc : blkif.rom_rdata <= 32'h93001000;
          16'h04cd : blkif.rom_rdata <= 32'h639a0000;
          16'h04ce : blkif.rom_rdata <= 32'h93801000;
          16'h04cf : blkif.rom_rdata <= 32'h93801000;
          16'h04d0 : blkif.rom_rdata <= 32'h93801000;
          16'h04d1 : blkif.rom_rdata <= 32'h93801000;
          16'h04d2 : blkif.rom_rdata <= 32'h93801000;
          16'h04d3 : blkif.rom_rdata <= 32'h93801000;
          16'h04d4 : blkif.rom_rdata <= 32'h930e3000;
          16'h04d5 : blkif.rom_rdata <= 32'h130e500e;
          16'h04d6 : blkif.rom_rdata <= 32'h6384d001;
          16'h04d7 : blkif.rom_rdata <= 32'h6f400041;
          16'h04d8 : blkif.rom_rdata <= 32'hb7000080;
          16'h04d9 : blkif.rom_rdata <= 32'h93804000;
          16'h04da : blkif.rom_rdata <= 32'h1301e001;
          16'h04db : blkif.rom_rdata <= 32'h23a02000;
          16'h04dc : blkif.rom_rdata <= 32'hb7000080;
          16'h04dd : blkif.rom_rdata <= 32'h93804000;
          16'h04de : blkif.rom_rdata <= 32'h1301b00b;
          16'h04df : blkif.rom_rdata <= 32'h23a02000;
          16'h04e0 : blkif.rom_rdata <= 32'h73100034;
          16'h04e1 : blkif.rom_rdata <= 32'h9360000f;
          16'h04e2 : blkif.rom_rdata <= 32'h1361f000;
          16'h04e3 : blkif.rom_rdata <= 32'h93611000;
          16'h04e4 : blkif.rom_rdata <= 32'h1362f00f;
          16'h04e5 : blkif.rom_rdata <= 32'hf3a10034;
          16'h04e6 : blkif.rom_rdata <= 32'h63043000;
          16'h04e7 : blkif.rom_rdata <= 32'h6f40003d;
          16'h04e8 : blkif.rom_rdata <= 32'h93611000;
          16'h04e9 : blkif.rom_rdata <= 32'hf3210034;
          16'h04ea : blkif.rom_rdata <= 32'h63841100;
          16'h04eb : blkif.rom_rdata <= 32'h6f40003c;
          16'h04ec : blkif.rom_rdata <= 32'hf3210134;
          16'h04ed : blkif.rom_rdata <= 32'h63841100;
          16'h04ee : blkif.rom_rdata <= 32'h6f40403b;
          16'h04ef : blkif.rom_rdata <= 32'h130e800e;
          16'h04f0 : blkif.rom_rdata <= 32'h6f008000;
          16'h04f1 : blkif.rom_rdata <= 32'h6f40803a;
          16'h04f2 : blkif.rom_rdata <= 32'hb7000080;
          16'h04f3 : blkif.rom_rdata <= 32'h93804000;
          16'h04f4 : blkif.rom_rdata <= 32'h1301900e;
          16'h04f5 : blkif.rom_rdata <= 32'h23a02000;
          16'h04f6 : blkif.rom_rdata <= 32'h93001000;
          16'h04f7 : blkif.rom_rdata <= 32'h6f004001;
          16'h04f8 : blkif.rom_rdata <= 32'h93801000;
          16'h04f9 : blkif.rom_rdata <= 32'h93801000;
          16'h04fa : blkif.rom_rdata <= 32'h93801000;
          16'h04fb : blkif.rom_rdata <= 32'h93801000;
          16'h04fc : blkif.rom_rdata <= 32'h93801000;
          16'h04fd : blkif.rom_rdata <= 32'h93801000;
          16'h04fe : blkif.rom_rdata <= 32'h930e3000;
          16'h04ff : blkif.rom_rdata <= 32'h130e900e;
          16'h0500 : blkif.rom_rdata <= 32'h6384d001;
          16'h0501 : blkif.rom_rdata <= 32'h6f408036;
          16'h0502 : blkif.rom_rdata <= 32'h130ea00e;
          16'h0503 : blkif.rom_rdata <= 32'h93000000;
          16'h0504 : blkif.rom_rdata <= 32'hef000001;
          16'h0505 : blkif.rom_rdata <= 32'h13000000;
          16'h0506 : blkif.rom_rdata <= 32'h13000000;
          16'h0507 : blkif.rom_rdata <= 32'h6f400035;
          16'h0508 : blkif.rom_rdata <= 32'h17010000;
          16'h0509 : blkif.rom_rdata <= 32'h130101ff;
          16'h050a : blkif.rom_rdata <= 32'h13014100;
          16'h050b : blkif.rom_rdata <= 32'h63041100;
          16'h050c : blkif.rom_rdata <= 32'h6f40c033;
          16'h050d : blkif.rom_rdata <= 32'hb7000080;
          16'h050e : blkif.rom_rdata <= 32'h93804000;
          16'h050f : blkif.rom_rdata <= 32'h1301b00e;
          16'h0510 : blkif.rom_rdata <= 32'h23a02000;
          16'h0511 : blkif.rom_rdata <= 32'h13011000;
          16'h0512 : blkif.rom_rdata <= 32'hef004001;
          16'h0513 : blkif.rom_rdata <= 32'h13011100;
          16'h0514 : blkif.rom_rdata <= 32'h13011100;
          16'h0515 : blkif.rom_rdata <= 32'h13011100;
          16'h0516 : blkif.rom_rdata <= 32'h13011100;
          16'h0517 : blkif.rom_rdata <= 32'h13011100;
          16'h0518 : blkif.rom_rdata <= 32'h13011100;
          16'h0519 : blkif.rom_rdata <= 32'h930e3000;
          16'h051a : blkif.rom_rdata <= 32'h130eb00e;
          16'h051b : blkif.rom_rdata <= 32'h6304d101;
          16'h051c : blkif.rom_rdata <= 32'h6f40c02f;
          16'h051d : blkif.rom_rdata <= 32'h130ec00e;
          16'h051e : blkif.rom_rdata <= 32'h930f0000;
          16'h051f : blkif.rom_rdata <= 32'h17010000;
          16'h0520 : blkif.rom_rdata <= 32'h13018101;
          16'h0521 : blkif.rom_rdata <= 32'he7090100;
          16'h0522 : blkif.rom_rdata <= 32'h13000000;
          16'h0523 : blkif.rom_rdata <= 32'h13000000;
          16'h0524 : blkif.rom_rdata <= 32'h6f40c02d;
          16'h0525 : blkif.rom_rdata <= 32'h97000000;
          16'h0526 : blkif.rom_rdata <= 32'h938000ff;
          16'h0527 : blkif.rom_rdata <= 32'h93804000;
          16'h0528 : blkif.rom_rdata <= 32'h63843001;
          16'h0529 : blkif.rom_rdata <= 32'h6f40802c;
          16'h052a : blkif.rom_rdata <= 32'h130ed00e;
          16'h052b : blkif.rom_rdata <= 32'h930f0000;
          16'h052c : blkif.rom_rdata <= 32'h97010000;
          16'h052d : blkif.rom_rdata <= 32'h93814101;
          16'h052e : blkif.rom_rdata <= 32'h67800100;
          16'h052f : blkif.rom_rdata <= 32'h13000000;
          16'h0530 : blkif.rom_rdata <= 32'h6f40c02a;
          16'h0531 : blkif.rom_rdata <= 32'h63840f00;
          16'h0532 : blkif.rom_rdata <= 32'h6f40402a;
          16'h0533 : blkif.rom_rdata <= 32'h130ee00e;
          16'h0534 : blkif.rom_rdata <= 32'h13020000;
          16'h0535 : blkif.rom_rdata <= 32'h17030000;
          16'h0536 : blkif.rom_rdata <= 32'h13034301;
          16'h0537 : blkif.rom_rdata <= 32'he7090300;
          16'h0538 : blkif.rom_rdata <= 32'h6304c001;
          16'h0539 : blkif.rom_rdata <= 32'h6f408028;
          16'h053a : blkif.rom_rdata <= 32'h13021200;
          16'h053b : blkif.rom_rdata <= 32'h93022000;
          16'h053c : blkif.rom_rdata <= 32'he31252fe;
          16'h053d : blkif.rom_rdata <= 32'h130ef00e;
          16'h053e : blkif.rom_rdata <= 32'h13020000;
          16'h053f : blkif.rom_rdata <= 32'h17030000;
          16'h0540 : blkif.rom_rdata <= 32'h13038301;
          16'h0541 : blkif.rom_rdata <= 32'h13000000;
          16'h0542 : blkif.rom_rdata <= 32'he7090300;
          16'h0543 : blkif.rom_rdata <= 32'h6304c001;
          16'h0544 : blkif.rom_rdata <= 32'h6f40c025;
          16'h0545 : blkif.rom_rdata <= 32'h13021200;
          16'h0546 : blkif.rom_rdata <= 32'h93022000;
          16'h0547 : blkif.rom_rdata <= 32'he31052fe;
          16'h0548 : blkif.rom_rdata <= 32'h130e000f;
          16'h0549 : blkif.rom_rdata <= 32'h13020000;
          16'h054a : blkif.rom_rdata <= 32'h17030000;
          16'h054b : blkif.rom_rdata <= 32'h1303c301;
          16'h054c : blkif.rom_rdata <= 32'h13000000;
          16'h054d : blkif.rom_rdata <= 32'h13000000;
          16'h054e : blkif.rom_rdata <= 32'he7090300;
          16'h054f : blkif.rom_rdata <= 32'h6304c001;
          16'h0550 : blkif.rom_rdata <= 32'h6f40c022;
          16'h0551 : blkif.rom_rdata <= 32'h13021200;
          16'h0552 : blkif.rom_rdata <= 32'h93022000;
          16'h0553 : blkif.rom_rdata <= 32'he31e52fc;
          16'h0554 : blkif.rom_rdata <= 32'hb7000080;
          16'h0555 : blkif.rom_rdata <= 32'h93804000;
          16'h0556 : blkif.rom_rdata <= 32'h1301100f;
          16'h0557 : blkif.rom_rdata <= 32'h23a02000;
          16'h0558 : blkif.rom_rdata <= 32'h93001000;
          16'h0559 : blkif.rom_rdata <= 32'h17010000;
          16'h055a : blkif.rom_rdata <= 32'h1301c101;
          16'h055b : blkif.rom_rdata <= 32'he709c1ff;
          16'h055c : blkif.rom_rdata <= 32'h93801000;
          16'h055d : blkif.rom_rdata <= 32'h93801000;
          16'h055e : blkif.rom_rdata <= 32'h93801000;
          16'h055f : blkif.rom_rdata <= 32'h93801000;
          16'h0560 : blkif.rom_rdata <= 32'h93801000;
          16'h0561 : blkif.rom_rdata <= 32'h93801000;
          16'h0562 : blkif.rom_rdata <= 32'h930e4000;
          16'h0563 : blkif.rom_rdata <= 32'h130e100f;
          16'h0564 : blkif.rom_rdata <= 32'h6384d001;
          16'h0565 : blkif.rom_rdata <= 32'h6f40801d;
          16'h0566 : blkif.rom_rdata <= 32'hb7000080;
          16'h0567 : blkif.rom_rdata <= 32'h93804000;
          16'h0568 : blkif.rom_rdata <= 32'h1301200f;
          16'h0569 : blkif.rom_rdata <= 32'h23a02000;
          16'h056a : blkif.rom_rdata <= 32'h97500000;
          16'h056b : blkif.rom_rdata <= 32'h938000c0;
          16'h056c : blkif.rom_rdata <= 32'h83810000;
          16'h056d : blkif.rom_rdata <= 32'h930ef0ff;
          16'h056e : blkif.rom_rdata <= 32'h130e200f;
          16'h056f : blkif.rom_rdata <= 32'h6384d101;
          16'h0570 : blkif.rom_rdata <= 32'h6f40c01a;
          16'h0571 : blkif.rom_rdata <= 32'hb7000080;
          16'h0572 : blkif.rom_rdata <= 32'h93804000;
          16'h0573 : blkif.rom_rdata <= 32'h1301500f;
          16'h0574 : blkif.rom_rdata <= 32'h23a02000;
          16'h0575 : blkif.rom_rdata <= 32'h97500000;
          16'h0576 : blkif.rom_rdata <= 32'h938040bd;
          16'h0577 : blkif.rom_rdata <= 32'h83813000;
          16'h0578 : blkif.rom_rdata <= 32'h930ef000;
          16'h0579 : blkif.rom_rdata <= 32'h130e500f;
          16'h057a : blkif.rom_rdata <= 32'h6384d101;
          16'h057b : blkif.rom_rdata <= 32'h6f400018;
          16'h057c : blkif.rom_rdata <= 32'hb7000080;
          16'h057d : blkif.rom_rdata <= 32'h93804000;
          16'h057e : blkif.rom_rdata <= 32'h1301600f;
          16'h057f : blkif.rom_rdata <= 32'h23a02000;
          16'h0580 : blkif.rom_rdata <= 32'h97500000;
          16'h0581 : blkif.rom_rdata <= 32'h9380b0ba;
          16'h0582 : blkif.rom_rdata <= 32'h8381d0ff;
          16'h0583 : blkif.rom_rdata <= 32'h930ef0ff;
          16'h0584 : blkif.rom_rdata <= 32'h130e600f;
          16'h0585 : blkif.rom_rdata <= 32'h6384d101;
          16'h0586 : blkif.rom_rdata <= 32'h6f404015;
          16'h0587 : blkif.rom_rdata <= 32'hb7000080;
          16'h0588 : blkif.rom_rdata <= 32'h93804000;
          16'h0589 : blkif.rom_rdata <= 32'h1301900f;
          16'h058a : blkif.rom_rdata <= 32'h23a02000;
          16'h058b : blkif.rom_rdata <= 32'h97500000;
          16'h058c : blkif.rom_rdata <= 32'h9380f0b7;
          16'h058d : blkif.rom_rdata <= 32'h83810000;
          16'h058e : blkif.rom_rdata <= 32'h930ef000;
          16'h058f : blkif.rom_rdata <= 32'h130e900f;
          16'h0590 : blkif.rom_rdata <= 32'h6384d101;
          16'h0591 : blkif.rom_rdata <= 32'h6f408012;
          16'h0592 : blkif.rom_rdata <= 32'hb7000080;
          16'h0593 : blkif.rom_rdata <= 32'h93804000;
          16'h0594 : blkif.rom_rdata <= 32'h1301a00f;
          16'h0595 : blkif.rom_rdata <= 32'h23a02000;
          16'h0596 : blkif.rom_rdata <= 32'h97500000;
          16'h0597 : blkif.rom_rdata <= 32'h938000b5;
          16'h0598 : blkif.rom_rdata <= 32'h938000fe;
          16'h0599 : blkif.rom_rdata <= 32'h83810002;
          16'h059a : blkif.rom_rdata <= 32'h930ef0ff;
          16'h059b : blkif.rom_rdata <= 32'h130ea00f;
          16'h059c : blkif.rom_rdata <= 32'h6384d101;
          16'h059d : blkif.rom_rdata <= 32'h6f40800f;
          16'h059e : blkif.rom_rdata <= 32'hb7000080;
          16'h059f : blkif.rom_rdata <= 32'h93804000;
          16'h05a0 : blkif.rom_rdata <= 32'h1301b00f;
          16'h05a1 : blkif.rom_rdata <= 32'h23a02000;
          16'h05a2 : blkif.rom_rdata <= 32'h97500000;
          16'h05a3 : blkif.rom_rdata <= 32'h938000b2;
          16'h05a4 : blkif.rom_rdata <= 32'h9380a0ff;
          16'h05a5 : blkif.rom_rdata <= 32'h83817000;
          16'h05a6 : blkif.rom_rdata <= 32'h930e0000;
          16'h05a7 : blkif.rom_rdata <= 32'h130eb00f;
          16'h05a8 : blkif.rom_rdata <= 32'h6384d101;
          16'h05a9 : blkif.rom_rdata <= 32'h6f40800c;
          16'h05aa : blkif.rom_rdata <= 32'h130ec00f;
          16'h05ab : blkif.rom_rdata <= 32'h13020000;
          16'h05ac : blkif.rom_rdata <= 32'h97500000;
          16'h05ad : blkif.rom_rdata <= 32'h938090af;
          16'h05ae : blkif.rom_rdata <= 32'h83811000;
          16'h05af : blkif.rom_rdata <= 32'h13830100;
          16'h05b0 : blkif.rom_rdata <= 32'h930e00ff;
          16'h05b1 : blkif.rom_rdata <= 32'h6304d301;
          16'h05b2 : blkif.rom_rdata <= 32'h6f40400a;
          16'h05b3 : blkif.rom_rdata <= 32'h13021200;
          16'h05b4 : blkif.rom_rdata <= 32'h93022000;
          16'h05b5 : blkif.rom_rdata <= 32'he31e52fc;
          16'h05b6 : blkif.rom_rdata <= 32'h130ee00f;
          16'h05b7 : blkif.rom_rdata <= 32'h13020000;
          16'h05b8 : blkif.rom_rdata <= 32'h97500000;
          16'h05b9 : blkif.rom_rdata <= 32'h938080ac;
          16'h05ba : blkif.rom_rdata <= 32'h83811000;
          16'h05bb : blkif.rom_rdata <= 32'h13000000;
          16'h05bc : blkif.rom_rdata <= 32'h13000000;
          16'h05bd : blkif.rom_rdata <= 32'h13830100;
          16'h05be : blkif.rom_rdata <= 32'h930e0000;
          16'h05bf : blkif.rom_rdata <= 32'h6304d301;
          16'h05c0 : blkif.rom_rdata <= 32'h6f40c006;
          16'h05c1 : blkif.rom_rdata <= 32'h13021200;
          16'h05c2 : blkif.rom_rdata <= 32'h93022000;
          16'h05c3 : blkif.rom_rdata <= 32'he31a52fc;
          16'h05c4 : blkif.rom_rdata <= 32'h130e0010;
          16'h05c5 : blkif.rom_rdata <= 32'h13020000;
          16'h05c6 : blkif.rom_rdata <= 32'h97500000;
          16'h05c7 : blkif.rom_rdata <= 32'h938020a9;
          16'h05c8 : blkif.rom_rdata <= 32'h13000000;
          16'h05c9 : blkif.rom_rdata <= 32'h83811000;
          16'h05ca : blkif.rom_rdata <= 32'h930ef000;
          16'h05cb : blkif.rom_rdata <= 32'h6384d101;
          16'h05cc : blkif.rom_rdata <= 32'h6f40c003;
          16'h05cd : blkif.rom_rdata <= 32'h13021200;
          16'h05ce : blkif.rom_rdata <= 32'h93022000;
          16'h05cf : blkif.rom_rdata <= 32'he31e52fc;
          16'h05d0 : blkif.rom_rdata <= 32'h130e1010;
          16'h05d1 : blkif.rom_rdata <= 32'h13020000;
          16'h05d2 : blkif.rom_rdata <= 32'h97500000;
          16'h05d3 : blkif.rom_rdata <= 32'h938000a6;
          16'h05d4 : blkif.rom_rdata <= 32'h13000000;
          16'h05d5 : blkif.rom_rdata <= 32'h13000000;
          16'h05d6 : blkif.rom_rdata <= 32'h83811000;
          16'h05d7 : blkif.rom_rdata <= 32'h930e0000;
          16'h05d8 : blkif.rom_rdata <= 32'h6384d101;
          16'h05d9 : blkif.rom_rdata <= 32'h6f408000;
          16'h05da : blkif.rom_rdata <= 32'h13021200;
          16'h05db : blkif.rom_rdata <= 32'h93022000;
          16'h05dc : blkif.rom_rdata <= 32'he31c52fc;
          16'h05dd : blkif.rom_rdata <= 32'hb7000080;
          16'h05de : blkif.rom_rdata <= 32'h93804000;
          16'h05df : blkif.rom_rdata <= 32'h13012010;
          16'h05e0 : blkif.rom_rdata <= 32'h23a02000;
          16'h05e1 : blkif.rom_rdata <= 32'h97510000;
          16'h05e2 : blkif.rom_rdata <= 32'h938141a2;
          16'h05e3 : blkif.rom_rdata <= 32'h03810100;
          16'h05e4 : blkif.rom_rdata <= 32'h13012000;
          16'h05e5 : blkif.rom_rdata <= 32'h930e2000;
          16'h05e6 : blkif.rom_rdata <= 32'h130e2010;
          16'h05e7 : blkif.rom_rdata <= 32'h6304d101;
          16'h05e8 : blkif.rom_rdata <= 32'h6f30d07c;
          16'h05e9 : blkif.rom_rdata <= 32'hb7000080;
          16'h05ea : blkif.rom_rdata <= 32'h93804000;
          16'h05eb : blkif.rom_rdata <= 32'h13013010;
          16'h05ec : blkif.rom_rdata <= 32'h23a02000;
          16'h05ed : blkif.rom_rdata <= 32'h97510000;
          16'h05ee : blkif.rom_rdata <= 32'h9381419f;
          16'h05ef : blkif.rom_rdata <= 32'h03810100;
          16'h05f0 : blkif.rom_rdata <= 32'h13000000;
          16'h05f1 : blkif.rom_rdata <= 32'h13012000;
          16'h05f2 : blkif.rom_rdata <= 32'h930e2000;
          16'h05f3 : blkif.rom_rdata <= 32'h130e3010;
          16'h05f4 : blkif.rom_rdata <= 32'h6304d101;
          16'h05f5 : blkif.rom_rdata <= 32'h6f309079;
          16'h05f6 : blkif.rom_rdata <= 32'hb7000080;
          16'h05f7 : blkif.rom_rdata <= 32'h93804000;
          16'h05f8 : blkif.rom_rdata <= 32'h13014010;
          16'h05f9 : blkif.rom_rdata <= 32'h23a02000;
          16'h05fa : blkif.rom_rdata <= 32'h97500000;
          16'h05fb : blkif.rom_rdata <= 32'h9380409c;
          16'h05fc : blkif.rom_rdata <= 32'h83c10000;
          16'h05fd : blkif.rom_rdata <= 32'h930ef00f;
          16'h05fe : blkif.rom_rdata <= 32'h130e4010;
          16'h05ff : blkif.rom_rdata <= 32'h6384d101;
          16'h0600 : blkif.rom_rdata <= 32'h6f30d076;
          16'h0601 : blkif.rom_rdata <= 32'hb7000080;
          16'h0602 : blkif.rom_rdata <= 32'h93804000;
          16'h0603 : blkif.rom_rdata <= 32'h13017010;
          16'h0604 : blkif.rom_rdata <= 32'h23a02000;
          16'h0605 : blkif.rom_rdata <= 32'h97500000;
          16'h0606 : blkif.rom_rdata <= 32'h93808099;
          16'h0607 : blkif.rom_rdata <= 32'h83c13000;
          16'h0608 : blkif.rom_rdata <= 32'h930ef000;
          16'h0609 : blkif.rom_rdata <= 32'h130e7010;
          16'h060a : blkif.rom_rdata <= 32'h6384d101;
          16'h060b : blkif.rom_rdata <= 32'h6f301074;
          16'h060c : blkif.rom_rdata <= 32'hb7000080;
          16'h060d : blkif.rom_rdata <= 32'h93804000;
          16'h060e : blkif.rom_rdata <= 32'h13018010;
          16'h060f : blkif.rom_rdata <= 32'h23a02000;
          16'h0610 : blkif.rom_rdata <= 32'h97500000;
          16'h0611 : blkif.rom_rdata <= 32'h9380f096;
          16'h0612 : blkif.rom_rdata <= 32'h83c1d0ff;
          16'h0613 : blkif.rom_rdata <= 32'h930ef00f;
          16'h0614 : blkif.rom_rdata <= 32'h130e8010;
          16'h0615 : blkif.rom_rdata <= 32'h6384d101;
          16'h0616 : blkif.rom_rdata <= 32'h6f305071;
          16'h0617 : blkif.rom_rdata <= 32'hb7000080;
          16'h0618 : blkif.rom_rdata <= 32'h93804000;
          16'h0619 : blkif.rom_rdata <= 32'h1301a010;
          16'h061a : blkif.rom_rdata <= 32'h23a02000;
          16'h061b : blkif.rom_rdata <= 32'h97500000;
          16'h061c : blkif.rom_rdata <= 32'h93803094;
          16'h061d : blkif.rom_rdata <= 32'h83c1f0ff;
          16'h061e : blkif.rom_rdata <= 32'h930e000f;
          16'h061f : blkif.rom_rdata <= 32'h130ea010;
          16'h0620 : blkif.rom_rdata <= 32'h6384d101;
          16'h0621 : blkif.rom_rdata <= 32'h6f30906e;
          16'h0622 : blkif.rom_rdata <= 32'hb7000080;
          16'h0623 : blkif.rom_rdata <= 32'h93804000;
          16'h0624 : blkif.rom_rdata <= 32'h1301c010;
          16'h0625 : blkif.rom_rdata <= 32'h23a02000;
          16'h0626 : blkif.rom_rdata <= 32'h97500000;
          16'h0627 : blkif.rom_rdata <= 32'h93804091;
          16'h0628 : blkif.rom_rdata <= 32'h938000fe;
          16'h0629 : blkif.rom_rdata <= 32'h83c10002;
          16'h062a : blkif.rom_rdata <= 32'h930ef00f;
          16'h062b : blkif.rom_rdata <= 32'h130ec010;
          16'h062c : blkif.rom_rdata <= 32'h6384d101;
          16'h062d : blkif.rom_rdata <= 32'h6f30906b;
          16'h062e : blkif.rom_rdata <= 32'hb7000080;
          16'h062f : blkif.rom_rdata <= 32'h93804000;
          16'h0630 : blkif.rom_rdata <= 32'h1301d010;
          16'h0631 : blkif.rom_rdata <= 32'h23a02000;
          16'h0632 : blkif.rom_rdata <= 32'h97500000;
          16'h0633 : blkif.rom_rdata <= 32'h9380408e;
          16'h0634 : blkif.rom_rdata <= 32'h9380a0ff;
          16'h0635 : blkif.rom_rdata <= 32'h83c17000;
          16'h0636 : blkif.rom_rdata <= 32'h930e0000;
          16'h0637 : blkif.rom_rdata <= 32'h130ed010;
          16'h0638 : blkif.rom_rdata <= 32'h6384d101;
          16'h0639 : blkif.rom_rdata <= 32'h6f309068;
          16'h063a : blkif.rom_rdata <= 32'h130ee010;
          16'h063b : blkif.rom_rdata <= 32'h13020000;
          16'h063c : blkif.rom_rdata <= 32'h97500000;
          16'h063d : blkif.rom_rdata <= 32'h9380d08b;
          16'h063e : blkif.rom_rdata <= 32'h83c11000;
          16'h063f : blkif.rom_rdata <= 32'h13830100;
          16'h0640 : blkif.rom_rdata <= 32'h930e000f;
          16'h0641 : blkif.rom_rdata <= 32'h6304d301;
          16'h0642 : blkif.rom_rdata <= 32'h6f305066;
          16'h0643 : blkif.rom_rdata <= 32'h13021200;
          16'h0644 : blkif.rom_rdata <= 32'h93022000;
          16'h0645 : blkif.rom_rdata <= 32'he31e52fc;
          16'h0646 : blkif.rom_rdata <= 32'h130e0011;
          16'h0647 : blkif.rom_rdata <= 32'h13020000;
          16'h0648 : blkif.rom_rdata <= 32'h97500000;
          16'h0649 : blkif.rom_rdata <= 32'h9380c088;
          16'h064a : blkif.rom_rdata <= 32'h83c11000;
          16'h064b : blkif.rom_rdata <= 32'h13000000;
          16'h064c : blkif.rom_rdata <= 32'h13000000;
          16'h064d : blkif.rom_rdata <= 32'h13830100;
          16'h064e : blkif.rom_rdata <= 32'h930e0000;
          16'h064f : blkif.rom_rdata <= 32'h6304d301;
          16'h0650 : blkif.rom_rdata <= 32'h6f30d062;
          16'h0651 : blkif.rom_rdata <= 32'h13021200;
          16'h0652 : blkif.rom_rdata <= 32'h93022000;
          16'h0653 : blkif.rom_rdata <= 32'he31a52fc;
          16'h0654 : blkif.rom_rdata <= 32'h130e1011;
          16'h0655 : blkif.rom_rdata <= 32'h13020000;
          16'h0656 : blkif.rom_rdata <= 32'h97500000;
          16'h0657 : blkif.rom_rdata <= 32'h93805085;
          16'h0658 : blkif.rom_rdata <= 32'h83c11000;
          16'h0659 : blkif.rom_rdata <= 32'h930e000f;
          16'h065a : blkif.rom_rdata <= 32'h6384d101;
          16'h065b : blkif.rom_rdata <= 32'h6f301060;
          16'h065c : blkif.rom_rdata <= 32'h13021200;
          16'h065d : blkif.rom_rdata <= 32'h93022000;
          16'h065e : blkif.rom_rdata <= 32'he31052fe;
          16'h065f : blkif.rom_rdata <= 32'h130e2011;
          16'h0660 : blkif.rom_rdata <= 32'h13020000;
          16'h0661 : blkif.rom_rdata <= 32'h97500000;
          16'h0662 : blkif.rom_rdata <= 32'h9380a082;
          16'h0663 : blkif.rom_rdata <= 32'h13000000;
          16'h0664 : blkif.rom_rdata <= 32'h83c11000;
          16'h0665 : blkif.rom_rdata <= 32'h930ef000;
          16'h0666 : blkif.rom_rdata <= 32'h6384d101;
          16'h0667 : blkif.rom_rdata <= 32'h6f30105d;
          16'h0668 : blkif.rom_rdata <= 32'h13021200;
          16'h0669 : blkif.rom_rdata <= 32'h93022000;
          16'h066a : blkif.rom_rdata <= 32'he31e52fc;
          16'h066b : blkif.rom_rdata <= 32'hb7000080;
          16'h066c : blkif.rom_rdata <= 32'h93804000;
          16'h066d : blkif.rom_rdata <= 32'h13014011;
          16'h066e : blkif.rom_rdata <= 32'h23a02000;
          16'h066f : blkif.rom_rdata <= 32'h97410000;
          16'h0670 : blkif.rom_rdata <= 32'h9381017f;
          16'h0671 : blkif.rom_rdata <= 32'h03c10100;
          16'h0672 : blkif.rom_rdata <= 32'h13012000;
          16'h0673 : blkif.rom_rdata <= 32'h930e2000;
          16'h0674 : blkif.rom_rdata <= 32'h130e4011;
          16'h0675 : blkif.rom_rdata <= 32'h6304d101;
          16'h0676 : blkif.rom_rdata <= 32'h6f305059;
          16'h0677 : blkif.rom_rdata <= 32'hb7000080;
          16'h0678 : blkif.rom_rdata <= 32'h93804000;
          16'h0679 : blkif.rom_rdata <= 32'h13015011;
          16'h067a : blkif.rom_rdata <= 32'h23a02000;
          16'h067b : blkif.rom_rdata <= 32'h97410000;
          16'h067c : blkif.rom_rdata <= 32'h9381017c;
          16'h067d : blkif.rom_rdata <= 32'h03c10100;
          16'h067e : blkif.rom_rdata <= 32'h13000000;
          16'h067f : blkif.rom_rdata <= 32'h13012000;
          16'h0680 : blkif.rom_rdata <= 32'h930e2000;
          16'h0681 : blkif.rom_rdata <= 32'h130e5011;
          16'h0682 : blkif.rom_rdata <= 32'h6304d101;
          16'h0683 : blkif.rom_rdata <= 32'h6f301056;
          16'h0684 : blkif.rom_rdata <= 32'hb7000080;
          16'h0685 : blkif.rom_rdata <= 32'h93804000;
          16'h0686 : blkif.rom_rdata <= 32'h13016011;
          16'h0687 : blkif.rom_rdata <= 32'h23a02000;
          16'h0688 : blkif.rom_rdata <= 32'h97400000;
          16'h0689 : blkif.rom_rdata <= 32'h93800079;
          16'h068a : blkif.rom_rdata <= 32'h83910000;
          16'h068b : blkif.rom_rdata <= 32'h930ef00f;
          16'h068c : blkif.rom_rdata <= 32'h130e6011;
          16'h068d : blkif.rom_rdata <= 32'h6384d101;
          16'h068e : blkif.rom_rdata <= 32'h6f305053;
          16'h068f : blkif.rom_rdata <= 32'hb7000080;
          16'h0690 : blkif.rom_rdata <= 32'h93804000;
          16'h0691 : blkif.rom_rdata <= 32'h13017011;
          16'h0692 : blkif.rom_rdata <= 32'h23a02000;
          16'h0693 : blkif.rom_rdata <= 32'h97400000;
          16'h0694 : blkif.rom_rdata <= 32'h93804076;
          16'h0695 : blkif.rom_rdata <= 32'h83912000;
          16'h0696 : blkif.rom_rdata <= 32'h930e00f0;
          16'h0697 : blkif.rom_rdata <= 32'h130e7011;
          16'h0698 : blkif.rom_rdata <= 32'h6384d101;
          16'h0699 : blkif.rom_rdata <= 32'h6f309050;
          16'h069a : blkif.rom_rdata <= 32'hb7000080;
          16'h069b : blkif.rom_rdata <= 32'h93804000;
          16'h069c : blkif.rom_rdata <= 32'h13019011;
          16'h069d : blkif.rom_rdata <= 32'h23a02000;
          16'h069e : blkif.rom_rdata <= 32'h97400000;
          16'h069f : blkif.rom_rdata <= 32'h93808073;
          16'h06a0 : blkif.rom_rdata <= 32'h83916000;
          16'h06a1 : blkif.rom_rdata <= 32'hb7feffff;
          16'h06a2 : blkif.rom_rdata <= 32'h938efe00;
          16'h06a3 : blkif.rom_rdata <= 32'h130e9011;
          16'h06a4 : blkif.rom_rdata <= 32'h6384d101;
          16'h06a5 : blkif.rom_rdata <= 32'h6f30904d;
          16'h06a6 : blkif.rom_rdata <= 32'hb7000080;
          16'h06a7 : blkif.rom_rdata <= 32'h93804000;
          16'h06a8 : blkif.rom_rdata <= 32'h1301a011;
          16'h06a9 : blkif.rom_rdata <= 32'h23a02000;
          16'h06aa : blkif.rom_rdata <= 32'h97400000;
          16'h06ab : blkif.rom_rdata <= 32'h9380e070;
          16'h06ac : blkif.rom_rdata <= 32'h8391a0ff;
          16'h06ad : blkif.rom_rdata <= 32'h930ef00f;
          16'h06ae : blkif.rom_rdata <= 32'h130ea011;
          16'h06af : blkif.rom_rdata <= 32'h6384d101;
          16'h06b0 : blkif.rom_rdata <= 32'h6f30d04a;
          16'h06b1 : blkif.rom_rdata <= 32'hb7000080;
          16'h06b2 : blkif.rom_rdata <= 32'h93804000;
          16'h06b3 : blkif.rom_rdata <= 32'h1301c011;
          16'h06b4 : blkif.rom_rdata <= 32'h23a02000;
          16'h06b5 : blkif.rom_rdata <= 32'h97400000;
          16'h06b6 : blkif.rom_rdata <= 32'h9380206e;
          16'h06b7 : blkif.rom_rdata <= 32'h8391e0ff;
          16'h06b8 : blkif.rom_rdata <= 32'hb71e0000;
          16'h06b9 : blkif.rom_rdata <= 32'h938e0eff;
          16'h06ba : blkif.rom_rdata <= 32'h130ec011;
          16'h06bb : blkif.rom_rdata <= 32'h6384d101;
          16'h06bc : blkif.rom_rdata <= 32'h6f30d047;
          16'h06bd : blkif.rom_rdata <= 32'hb7000080;
          16'h06be : blkif.rom_rdata <= 32'h93804000;
          16'h06bf : blkif.rom_rdata <= 32'h1301d011;
          16'h06c0 : blkif.rom_rdata <= 32'h23a02000;
          16'h06c1 : blkif.rom_rdata <= 32'h97400000;
          16'h06c2 : blkif.rom_rdata <= 32'h9380206b;
          16'h06c3 : blkif.rom_rdata <= 32'h83910000;
          16'h06c4 : blkif.rom_rdata <= 32'hb7feffff;
          16'h06c5 : blkif.rom_rdata <= 32'h938efe00;
          16'h06c6 : blkif.rom_rdata <= 32'h130ed011;
          16'h06c7 : blkif.rom_rdata <= 32'h6384d101;
          16'h06c8 : blkif.rom_rdata <= 32'h6f30d044;
          16'h06c9 : blkif.rom_rdata <= 32'hb7000080;
          16'h06ca : blkif.rom_rdata <= 32'h93804000;
          16'h06cb : blkif.rom_rdata <= 32'h1301e011;
          16'h06cc : blkif.rom_rdata <= 32'h23a02000;
          16'h06cd : blkif.rom_rdata <= 32'h97400000;
          16'h06ce : blkif.rom_rdata <= 32'h9380c067;
          16'h06cf : blkif.rom_rdata <= 32'h938000fe;
          16'h06d0 : blkif.rom_rdata <= 32'h83910002;
          16'h06d1 : blkif.rom_rdata <= 32'h930ef00f;
          16'h06d2 : blkif.rom_rdata <= 32'h130ee011;
          16'h06d3 : blkif.rom_rdata <= 32'h6384d101;
          16'h06d4 : blkif.rom_rdata <= 32'h6f30d041;
          16'h06d5 : blkif.rom_rdata <= 32'hb7000080;
          16'h06d6 : blkif.rom_rdata <= 32'h93804000;
          16'h06d7 : blkif.rom_rdata <= 32'h1301f011;
          16'h06d8 : blkif.rom_rdata <= 32'h23a02000;
          16'h06d9 : blkif.rom_rdata <= 32'h97400000;
          16'h06da : blkif.rom_rdata <= 32'h9380c064;
          16'h06db : blkif.rom_rdata <= 32'h9380b0ff;
          16'h06dc : blkif.rom_rdata <= 32'h83917000;
          16'h06dd : blkif.rom_rdata <= 32'h930e00f0;
          16'h06de : blkif.rom_rdata <= 32'h130ef011;
          16'h06df : blkif.rom_rdata <= 32'h6384d101;
          16'h06e0 : blkif.rom_rdata <= 32'h6f30d03e;
          16'h06e1 : blkif.rom_rdata <= 32'h130e0012;
          16'h06e2 : blkif.rom_rdata <= 32'h13020000;
          16'h06e3 : blkif.rom_rdata <= 32'h97400000;
          16'h06e4 : blkif.rom_rdata <= 32'h93806062;
          16'h06e5 : blkif.rom_rdata <= 32'h83912000;
          16'h06e6 : blkif.rom_rdata <= 32'h13830100;
          16'h06e7 : blkif.rom_rdata <= 32'hb71e0000;
          16'h06e8 : blkif.rom_rdata <= 32'h938e0eff;
          16'h06e9 : blkif.rom_rdata <= 32'h6304d301;
          16'h06ea : blkif.rom_rdata <= 32'h6f30503c;
          16'h06eb : blkif.rom_rdata <= 32'h13021200;
          16'h06ec : blkif.rom_rdata <= 32'h93022000;
          16'h06ed : blkif.rom_rdata <= 32'he31c52fc;
          16'h06ee : blkif.rom_rdata <= 32'h130e2012;
          16'h06ef : blkif.rom_rdata <= 32'h13020000;
          16'h06f0 : blkif.rom_rdata <= 32'h97400000;
          16'h06f1 : blkif.rom_rdata <= 32'h9380005f;
          16'h06f2 : blkif.rom_rdata <= 32'h83912000;
          16'h06f3 : blkif.rom_rdata <= 32'h13000000;
          16'h06f4 : blkif.rom_rdata <= 32'h13000000;
          16'h06f5 : blkif.rom_rdata <= 32'h13830100;
          16'h06f6 : blkif.rom_rdata <= 32'h930e00f0;
          16'h06f7 : blkif.rom_rdata <= 32'h6304d301;
          16'h06f8 : blkif.rom_rdata <= 32'h6f30d038;
          16'h06f9 : blkif.rom_rdata <= 32'h13021200;
          16'h06fa : blkif.rom_rdata <= 32'h93022000;
          16'h06fb : blkif.rom_rdata <= 32'he31a52fc;
          16'h06fc : blkif.rom_rdata <= 32'h130e4012;
          16'h06fd : blkif.rom_rdata <= 32'h13020000;
          16'h06fe : blkif.rom_rdata <= 32'h97400000;
          16'h06ff : blkif.rom_rdata <= 32'h9380c05b;
          16'h0700 : blkif.rom_rdata <= 32'h13000000;
          16'h0701 : blkif.rom_rdata <= 32'h83912000;
          16'h0702 : blkif.rom_rdata <= 32'hb7feffff;
          16'h0703 : blkif.rom_rdata <= 32'h938efe00;
          16'h0704 : blkif.rom_rdata <= 32'h6384d101;
          16'h0705 : blkif.rom_rdata <= 32'h6f309035;
          16'h0706 : blkif.rom_rdata <= 32'h13021200;
          16'h0707 : blkif.rom_rdata <= 32'h93022000;
          16'h0708 : blkif.rom_rdata <= 32'he31c52fc;
          16'h0709 : blkif.rom_rdata <= 32'h130e5012;
          16'h070a : blkif.rom_rdata <= 32'h13020000;
          16'h070b : blkif.rom_rdata <= 32'h97400000;
          16'h070c : blkif.rom_rdata <= 32'h93804058;
          16'h070d : blkif.rom_rdata <= 32'h13000000;
          16'h070e : blkif.rom_rdata <= 32'h13000000;
          16'h070f : blkif.rom_rdata <= 32'h83912000;
          16'h0710 : blkif.rom_rdata <= 32'h930e00f0;
          16'h0711 : blkif.rom_rdata <= 32'h6384d101;
          16'h0712 : blkif.rom_rdata <= 32'h6f305032;
          16'h0713 : blkif.rom_rdata <= 32'h13021200;
          16'h0714 : blkif.rom_rdata <= 32'h93022000;
          16'h0715 : blkif.rom_rdata <= 32'he31c52fc;
          16'h0716 : blkif.rom_rdata <= 32'hb7000080;
          16'h0717 : blkif.rom_rdata <= 32'h93804000;
          16'h0718 : blkif.rom_rdata <= 32'h13016012;
          16'h0719 : blkif.rom_rdata <= 32'h23a02000;
          16'h071a : blkif.rom_rdata <= 32'h97410000;
          16'h071b : blkif.rom_rdata <= 32'h93818154;
          16'h071c : blkif.rom_rdata <= 32'h03910100;
          16'h071d : blkif.rom_rdata <= 32'h13012000;
          16'h071e : blkif.rom_rdata <= 32'h930e2000;
          16'h071f : blkif.rom_rdata <= 32'h130e6012;
          16'h0720 : blkif.rom_rdata <= 32'h6304d101;
          16'h0721 : blkif.rom_rdata <= 32'h6f30902e;
          16'h0722 : blkif.rom_rdata <= 32'hb7000080;
          16'h0723 : blkif.rom_rdata <= 32'h93804000;
          16'h0724 : blkif.rom_rdata <= 32'h13017012;
          16'h0725 : blkif.rom_rdata <= 32'h23a02000;
          16'h0726 : blkif.rom_rdata <= 32'h97410000;
          16'h0727 : blkif.rom_rdata <= 32'h93818151;
          16'h0728 : blkif.rom_rdata <= 32'h03910100;
          16'h0729 : blkif.rom_rdata <= 32'h13000000;
          16'h072a : blkif.rom_rdata <= 32'h13012000;
          16'h072b : blkif.rom_rdata <= 32'h930e2000;
          16'h072c : blkif.rom_rdata <= 32'h130e7012;
          16'h072d : blkif.rom_rdata <= 32'h6304d101;
          16'h072e : blkif.rom_rdata <= 32'h6f30502b;
          16'h072f : blkif.rom_rdata <= 32'hb7000080;
          16'h0730 : blkif.rom_rdata <= 32'h93804000;
          16'h0731 : blkif.rom_rdata <= 32'h13018012;
          16'h0732 : blkif.rom_rdata <= 32'h23a02000;
          16'h0733 : blkif.rom_rdata <= 32'h97400000;
          16'h0734 : blkif.rom_rdata <= 32'h9380c04e;
          16'h0735 : blkif.rom_rdata <= 32'h83d10000;
          16'h0736 : blkif.rom_rdata <= 32'h930ef00f;
          16'h0737 : blkif.rom_rdata <= 32'h130e8012;
          16'h0738 : blkif.rom_rdata <= 32'h6384d101;
          16'h0739 : blkif.rom_rdata <= 32'h6f309028;
          16'h073a : blkif.rom_rdata <= 32'hb7000080;
          16'h073b : blkif.rom_rdata <= 32'h93804000;
          16'h073c : blkif.rom_rdata <= 32'h13019012;
          16'h073d : blkif.rom_rdata <= 32'h23a02000;
          16'h073e : blkif.rom_rdata <= 32'h97400000;
          16'h073f : blkif.rom_rdata <= 32'h9380004c;
          16'h0740 : blkif.rom_rdata <= 32'h83d12000;
          16'h0741 : blkif.rom_rdata <= 32'hb70e0100;
          16'h0742 : blkif.rom_rdata <= 32'h938e0ef0;
          16'h0743 : blkif.rom_rdata <= 32'h130e9012;
          16'h0744 : blkif.rom_rdata <= 32'h6384d101;
          16'h0745 : blkif.rom_rdata <= 32'h6f309025;
          16'h0746 : blkif.rom_rdata <= 32'hb7000080;
          16'h0747 : blkif.rom_rdata <= 32'h93804000;
          16'h0748 : blkif.rom_rdata <= 32'h1301b012;
          16'h0749 : blkif.rom_rdata <= 32'h23a02000;
          16'h074a : blkif.rom_rdata <= 32'h97400000;
          16'h074b : blkif.rom_rdata <= 32'h93800049;
          16'h074c : blkif.rom_rdata <= 32'h83d16000;
          16'h074d : blkif.rom_rdata <= 32'hb7fe0000;
          16'h074e : blkif.rom_rdata <= 32'h938efe00;
          16'h074f : blkif.rom_rdata <= 32'h130eb012;
          16'h0750 : blkif.rom_rdata <= 32'h6384d101;
          16'h0751 : blkif.rom_rdata <= 32'h6f309022;
          16'h0752 : blkif.rom_rdata <= 32'hb7000080;
          16'h0753 : blkif.rom_rdata <= 32'h93804000;
          16'h0754 : blkif.rom_rdata <= 32'h1301c012;
          16'h0755 : blkif.rom_rdata <= 32'h23a02000;
          16'h0756 : blkif.rom_rdata <= 32'h97400000;
          16'h0757 : blkif.rom_rdata <= 32'h93806046;
          16'h0758 : blkif.rom_rdata <= 32'h83d1a0ff;
          16'h0759 : blkif.rom_rdata <= 32'h930ef00f;
          16'h075a : blkif.rom_rdata <= 32'h130ec012;
          16'h075b : blkif.rom_rdata <= 32'h6384d101;
          16'h075c : blkif.rom_rdata <= 32'h6f30d01f;
          16'h075d : blkif.rom_rdata <= 32'hb7000080;
          16'h075e : blkif.rom_rdata <= 32'h93804000;
          16'h075f : blkif.rom_rdata <= 32'h1301d012;
          16'h0760 : blkif.rom_rdata <= 32'h23a02000;
          16'h0761 : blkif.rom_rdata <= 32'h97400000;
          16'h0762 : blkif.rom_rdata <= 32'h9380a043;
          16'h0763 : blkif.rom_rdata <= 32'h83d1c0ff;
          16'h0764 : blkif.rom_rdata <= 32'hb70e0100;
          16'h0765 : blkif.rom_rdata <= 32'h938e0ef0;
          16'h0766 : blkif.rom_rdata <= 32'h130ed012;
          16'h0767 : blkif.rom_rdata <= 32'h6384d101;
          16'h0768 : blkif.rom_rdata <= 32'h6f30d01c;
          16'h0769 : blkif.rom_rdata <= 32'hb7000080;
          16'h076a : blkif.rom_rdata <= 32'h93804000;
          16'h076b : blkif.rom_rdata <= 32'h1301f012;
          16'h076c : blkif.rom_rdata <= 32'h23a02000;
          16'h076d : blkif.rom_rdata <= 32'h97400000;
          16'h076e : blkif.rom_rdata <= 32'h9380a040;
          16'h076f : blkif.rom_rdata <= 32'h83d10000;
          16'h0770 : blkif.rom_rdata <= 32'hb7fe0000;
          16'h0771 : blkif.rom_rdata <= 32'h938efe00;
          16'h0772 : blkif.rom_rdata <= 32'h130ef012;
          16'h0773 : blkif.rom_rdata <= 32'h6384d101;
          16'h0774 : blkif.rom_rdata <= 32'h6f30d019;
          16'h0775 : blkif.rom_rdata <= 32'hb7000080;
          16'h0776 : blkif.rom_rdata <= 32'h93804000;
          16'h0777 : blkif.rom_rdata <= 32'h13010013;
          16'h0778 : blkif.rom_rdata <= 32'h23a02000;
          16'h0779 : blkif.rom_rdata <= 32'h97400000;
          16'h077a : blkif.rom_rdata <= 32'h9380403d;
          16'h077b : blkif.rom_rdata <= 32'h938000fe;
          16'h077c : blkif.rom_rdata <= 32'h83d10002;
          16'h077d : blkif.rom_rdata <= 32'h930ef00f;
          16'h077e : blkif.rom_rdata <= 32'h130e0013;
          16'h077f : blkif.rom_rdata <= 32'h6384d101;
          16'h0780 : blkif.rom_rdata <= 32'h6f30d016;
          16'h0781 : blkif.rom_rdata <= 32'hb7000080;
          16'h0782 : blkif.rom_rdata <= 32'h93804000;
          16'h0783 : blkif.rom_rdata <= 32'h13011013;
          16'h0784 : blkif.rom_rdata <= 32'h23a02000;
          16'h0785 : blkif.rom_rdata <= 32'h97400000;
          16'h0786 : blkif.rom_rdata <= 32'h9380403a;
          16'h0787 : blkif.rom_rdata <= 32'h9380b0ff;
          16'h0788 : blkif.rom_rdata <= 32'h83d17000;
          16'h0789 : blkif.rom_rdata <= 32'hb70e0100;
          16'h078a : blkif.rom_rdata <= 32'h938e0ef0;
          16'h078b : blkif.rom_rdata <= 32'h130e1013;
          16'h078c : blkif.rom_rdata <= 32'h6384d101;
          16'h078d : blkif.rom_rdata <= 32'h6f309013;
          16'h078e : blkif.rom_rdata <= 32'h130e2013;
          16'h078f : blkif.rom_rdata <= 32'h13020000;
          16'h0790 : blkif.rom_rdata <= 32'h97400000;
          16'h0791 : blkif.rom_rdata <= 32'h9380a037;
          16'h0792 : blkif.rom_rdata <= 32'h83d12000;
          16'h0793 : blkif.rom_rdata <= 32'h13830100;
          16'h0794 : blkif.rom_rdata <= 32'hb71e0000;
          16'h0795 : blkif.rom_rdata <= 32'h938e0eff;
          16'h0796 : blkif.rom_rdata <= 32'h6304d301;
          16'h0797 : blkif.rom_rdata <= 32'h6f301011;
          16'h0798 : blkif.rom_rdata <= 32'h13021200;
          16'h0799 : blkif.rom_rdata <= 32'h93022000;
          16'h079a : blkif.rom_rdata <= 32'he31c52fc;
          16'h079b : blkif.rom_rdata <= 32'h130e4013;
          16'h079c : blkif.rom_rdata <= 32'h13020000;
          16'h079d : blkif.rom_rdata <= 32'h97400000;
          16'h079e : blkif.rom_rdata <= 32'h93804034;
          16'h079f : blkif.rom_rdata <= 32'h83d12000;
          16'h07a0 : blkif.rom_rdata <= 32'h13000000;
          16'h07a1 : blkif.rom_rdata <= 32'h13000000;
          16'h07a2 : blkif.rom_rdata <= 32'h13830100;
          16'h07a3 : blkif.rom_rdata <= 32'hb70e0100;
          16'h07a4 : blkif.rom_rdata <= 32'h938e0ef0;
          16'h07a5 : blkif.rom_rdata <= 32'h6304d301;
          16'h07a6 : blkif.rom_rdata <= 32'h6f30500d;
          16'h07a7 : blkif.rom_rdata <= 32'h13021200;
          16'h07a8 : blkif.rom_rdata <= 32'h93022000;
          16'h07a9 : blkif.rom_rdata <= 32'he31852fc;
          16'h07aa : blkif.rom_rdata <= 32'h130e5013;
          16'h07ab : blkif.rom_rdata <= 32'h13020000;
          16'h07ac : blkif.rom_rdata <= 32'h97400000;
          16'h07ad : blkif.rom_rdata <= 32'h9380a030;
          16'h07ae : blkif.rom_rdata <= 32'h83d12000;
          16'h07af : blkif.rom_rdata <= 32'hb71e0000;
          16'h07b0 : blkif.rom_rdata <= 32'h938e0eff;
          16'h07b1 : blkif.rom_rdata <= 32'h6384d101;
          16'h07b2 : blkif.rom_rdata <= 32'h6f30500a;
          16'h07b3 : blkif.rom_rdata <= 32'h13021200;
          16'h07b4 : blkif.rom_rdata <= 32'h93022000;
          16'h07b5 : blkif.rom_rdata <= 32'he31e52fc;
          16'h07b6 : blkif.rom_rdata <= 32'h130e6013;
          16'h07b7 : blkif.rom_rdata <= 32'h13020000;
          16'h07b8 : blkif.rom_rdata <= 32'h97400000;
          16'h07b9 : blkif.rom_rdata <= 32'h9380c02d;
          16'h07ba : blkif.rom_rdata <= 32'h13000000;
          16'h07bb : blkif.rom_rdata <= 32'h83d12000;
          16'h07bc : blkif.rom_rdata <= 32'hb7fe0000;
          16'h07bd : blkif.rom_rdata <= 32'h938efe00;
          16'h07be : blkif.rom_rdata <= 32'h6384d101;
          16'h07bf : blkif.rom_rdata <= 32'h6f301007;
          16'h07c0 : blkif.rom_rdata <= 32'h13021200;
          16'h07c1 : blkif.rom_rdata <= 32'h93022000;
          16'h07c2 : blkif.rom_rdata <= 32'he31c52fc;
          16'h07c3 : blkif.rom_rdata <= 32'h130e7013;
          16'h07c4 : blkif.rom_rdata <= 32'h13020000;
          16'h07c5 : blkif.rom_rdata <= 32'h97400000;
          16'h07c6 : blkif.rom_rdata <= 32'h9380402a;
          16'h07c7 : blkif.rom_rdata <= 32'h13000000;
          16'h07c8 : blkif.rom_rdata <= 32'h13000000;
          16'h07c9 : blkif.rom_rdata <= 32'h83d12000;
          16'h07ca : blkif.rom_rdata <= 32'hb70e0100;
          16'h07cb : blkif.rom_rdata <= 32'h938e0ef0;
          16'h07cc : blkif.rom_rdata <= 32'h6384d101;
          16'h07cd : blkif.rom_rdata <= 32'h6f309003;
          16'h07ce : blkif.rom_rdata <= 32'h13021200;
          16'h07cf : blkif.rom_rdata <= 32'h93022000;
          16'h07d0 : blkif.rom_rdata <= 32'he31a52fc;
          16'h07d1 : blkif.rom_rdata <= 32'hb7000080;
          16'h07d2 : blkif.rom_rdata <= 32'h93804000;
          16'h07d3 : blkif.rom_rdata <= 32'h13018013;
          16'h07d4 : blkif.rom_rdata <= 32'h23a02000;
          16'h07d5 : blkif.rom_rdata <= 32'h97410000;
          16'h07d6 : blkif.rom_rdata <= 32'h93814126;
          16'h07d7 : blkif.rom_rdata <= 32'h03d10100;
          16'h07d8 : blkif.rom_rdata <= 32'h13012000;
          16'h07d9 : blkif.rom_rdata <= 32'h930e2000;
          16'h07da : blkif.rom_rdata <= 32'h130e8013;
          16'h07db : blkif.rom_rdata <= 32'h6304d101;
          16'h07dc : blkif.rom_rdata <= 32'h6f30c07f;
          16'h07dd : blkif.rom_rdata <= 32'hb7000080;
          16'h07de : blkif.rom_rdata <= 32'h93804000;
          16'h07df : blkif.rom_rdata <= 32'h13019013;
          16'h07e0 : blkif.rom_rdata <= 32'h23a02000;
          16'h07e1 : blkif.rom_rdata <= 32'h97410000;
          16'h07e2 : blkif.rom_rdata <= 32'h93814123;
          16'h07e3 : blkif.rom_rdata <= 32'h03d10100;
          16'h07e4 : blkif.rom_rdata <= 32'h13000000;
          16'h07e5 : blkif.rom_rdata <= 32'h13012000;
          16'h07e6 : blkif.rom_rdata <= 32'h930e2000;
          16'h07e7 : blkif.rom_rdata <= 32'h130e9013;
          16'h07e8 : blkif.rom_rdata <= 32'h6304d101;
          16'h07e9 : blkif.rom_rdata <= 32'h6f30807c;
          16'h07ea : blkif.rom_rdata <= 32'hb7000080;
          16'h07eb : blkif.rom_rdata <= 32'h93804000;
          16'h07ec : blkif.rom_rdata <= 32'h1301a013;
          16'h07ed : blkif.rom_rdata <= 32'h23a02000;
          16'h07ee : blkif.rom_rdata <= 32'hb7000000;
          16'h07ef : blkif.rom_rdata <= 32'h930e0000;
          16'h07f0 : blkif.rom_rdata <= 32'h130ea013;
          16'h07f1 : blkif.rom_rdata <= 32'h6384d001;
          16'h07f2 : blkif.rom_rdata <= 32'h6f30407a;
          16'h07f3 : blkif.rom_rdata <= 32'hb7000080;
          16'h07f4 : blkif.rom_rdata <= 32'h93804000;
          16'h07f5 : blkif.rom_rdata <= 32'h1301b013;
          16'h07f6 : blkif.rom_rdata <= 32'h23a02000;
          16'h07f7 : blkif.rom_rdata <= 32'hb7f0ffff;
          16'h07f8 : blkif.rom_rdata <= 32'h93d01040;
          16'h07f9 : blkif.rom_rdata <= 32'h930e0080;
          16'h07fa : blkif.rom_rdata <= 32'h130eb013;
          16'h07fb : blkif.rom_rdata <= 32'h6384d001;
          16'h07fc : blkif.rom_rdata <= 32'h6f30c077;
          16'h07fd : blkif.rom_rdata <= 32'hb7000080;
          16'h07fe : blkif.rom_rdata <= 32'h93804000;
          16'h07ff : blkif.rom_rdata <= 32'h1301c013;
          16'h0800 : blkif.rom_rdata <= 32'h23a02000;
          16'h0801 : blkif.rom_rdata <= 32'hb7f0ff7f;
          16'h0802 : blkif.rom_rdata <= 32'h93d04041;
          16'h0803 : blkif.rom_rdata <= 32'h930ef07f;
          16'h0804 : blkif.rom_rdata <= 32'h130ec013;
          16'h0805 : blkif.rom_rdata <= 32'h6384d001;
          16'h0806 : blkif.rom_rdata <= 32'h6f304075;
          16'h0807 : blkif.rom_rdata <= 32'hb7000080;
          16'h0808 : blkif.rom_rdata <= 32'h93804000;
          16'h0809 : blkif.rom_rdata <= 32'h1301d013;
          16'h080a : blkif.rom_rdata <= 32'h23a02000;
          16'h080b : blkif.rom_rdata <= 32'hb7000080;
          16'h080c : blkif.rom_rdata <= 32'h93d04041;
          16'h080d : blkif.rom_rdata <= 32'h930e0080;
          16'h080e : blkif.rom_rdata <= 32'h130ed013;
          16'h080f : blkif.rom_rdata <= 32'h6384d001;
          16'h0810 : blkif.rom_rdata <= 32'h6f30c072;
          16'h0811 : blkif.rom_rdata <= 32'hb7000080;
          16'h0812 : blkif.rom_rdata <= 32'h93804000;
          16'h0813 : blkif.rom_rdata <= 32'h1301e013;
          16'h0814 : blkif.rom_rdata <= 32'h23a02000;
          16'h0815 : blkif.rom_rdata <= 32'h37000080;
          16'h0816 : blkif.rom_rdata <= 32'h930e0000;
          16'h0817 : blkif.rom_rdata <= 32'h130ee013;
          16'h0818 : blkif.rom_rdata <= 32'h6304d001;
          16'h0819 : blkif.rom_rdata <= 32'h6f308070;
          16'h081a : blkif.rom_rdata <= 32'hb7000080;
          16'h081b : blkif.rom_rdata <= 32'h93804000;
          16'h081c : blkif.rom_rdata <= 32'h1301f013;
          16'h081d : blkif.rom_rdata <= 32'h23a02000;
          16'h081e : blkif.rom_rdata <= 32'h97400000;
          16'h081f : blkif.rom_rdata <= 32'h93808014;
          16'h0820 : blkif.rom_rdata <= 32'h83a10000;
          16'h0821 : blkif.rom_rdata <= 32'hb70eff00;
          16'h0822 : blkif.rom_rdata <= 32'h938efe0f;
          16'h0823 : blkif.rom_rdata <= 32'h130ef013;
          16'h0824 : blkif.rom_rdata <= 32'h6384d101;
          16'h0825 : blkif.rom_rdata <= 32'h6f30806d;
          16'h0826 : blkif.rom_rdata <= 32'hb7000080;
          16'h0827 : blkif.rom_rdata <= 32'h93804000;
          16'h0828 : blkif.rom_rdata <= 32'h13012014;
          16'h0829 : blkif.rom_rdata <= 32'h23a02000;
          16'h082a : blkif.rom_rdata <= 32'h97400000;
          16'h082b : blkif.rom_rdata <= 32'h93808011;
          16'h082c : blkif.rom_rdata <= 32'h83a1c000;
          16'h082d : blkif.rom_rdata <= 32'hb7fe0ff0;
          16'h082e : blkif.rom_rdata <= 32'h938efe00;
          16'h082f : blkif.rom_rdata <= 32'h130e2014;
          16'h0830 : blkif.rom_rdata <= 32'h6384d101;
          16'h0831 : blkif.rom_rdata <= 32'h6f30806a;
          16'h0832 : blkif.rom_rdata <= 32'hb7000080;
          16'h0833 : blkif.rom_rdata <= 32'h93804000;
          16'h0834 : blkif.rom_rdata <= 32'h13014014;
          16'h0835 : blkif.rom_rdata <= 32'h23a02000;
          16'h0836 : blkif.rom_rdata <= 32'h97400000;
          16'h0837 : blkif.rom_rdata <= 32'h9380400f;
          16'h0838 : blkif.rom_rdata <= 32'h83a180ff;
          16'h0839 : blkif.rom_rdata <= 32'hb70e01ff;
          16'h083a : blkif.rom_rdata <= 32'h938e0ef0;
          16'h083b : blkif.rom_rdata <= 32'h130e4014;
          16'h083c : blkif.rom_rdata <= 32'h6384d101;
          16'h083d : blkif.rom_rdata <= 32'h6f308067;
          16'h083e : blkif.rom_rdata <= 32'hb7000080;
          16'h083f : blkif.rom_rdata <= 32'h93804000;
          16'h0840 : blkif.rom_rdata <= 32'h13016014;
          16'h0841 : blkif.rom_rdata <= 32'h23a02000;
          16'h0842 : blkif.rom_rdata <= 32'h97400000;
          16'h0843 : blkif.rom_rdata <= 32'h9380400c;
          16'h0844 : blkif.rom_rdata <= 32'h83a10000;
          16'h0845 : blkif.rom_rdata <= 32'hb7fe0ff0;
          16'h0846 : blkif.rom_rdata <= 32'h938efe00;
          16'h0847 : blkif.rom_rdata <= 32'h130e6014;
          16'h0848 : blkif.rom_rdata <= 32'h6384d101;
          16'h0849 : blkif.rom_rdata <= 32'h6f308064;
          16'h084a : blkif.rom_rdata <= 32'hb7000080;
          16'h084b : blkif.rom_rdata <= 32'h93804000;
          16'h084c : blkif.rom_rdata <= 32'h13017014;
          16'h084d : blkif.rom_rdata <= 32'h23a02000;
          16'h084e : blkif.rom_rdata <= 32'h97400000;
          16'h084f : blkif.rom_rdata <= 32'h93808008;
          16'h0850 : blkif.rom_rdata <= 32'h938000fe;
          16'h0851 : blkif.rom_rdata <= 32'h83a10002;
          16'h0852 : blkif.rom_rdata <= 32'hb70eff00;
          16'h0853 : blkif.rom_rdata <= 32'h938efe0f;
          16'h0854 : blkif.rom_rdata <= 32'h130e7014;
          16'h0855 : blkif.rom_rdata <= 32'h6384d101;
          16'h0856 : blkif.rom_rdata <= 32'h6f304061;
          16'h0857 : blkif.rom_rdata <= 32'hb7000080;
          16'h0858 : blkif.rom_rdata <= 32'h93804000;
          16'h0859 : blkif.rom_rdata <= 32'h13018014;
          16'h085a : blkif.rom_rdata <= 32'h23a02000;
          16'h085b : blkif.rom_rdata <= 32'h97400000;
          16'h085c : blkif.rom_rdata <= 32'h93804005;
          16'h085d : blkif.rom_rdata <= 32'h9380d0ff;
          16'h085e : blkif.rom_rdata <= 32'h83a17000;
          16'h085f : blkif.rom_rdata <= 32'hb70e01ff;
          16'h0860 : blkif.rom_rdata <= 32'h938e0ef0;
          16'h0861 : blkif.rom_rdata <= 32'h130e8014;
          16'h0862 : blkif.rom_rdata <= 32'h6384d101;
          16'h0863 : blkif.rom_rdata <= 32'h6f30005e;
          16'h0864 : blkif.rom_rdata <= 32'h130e9014;
          16'h0865 : blkif.rom_rdata <= 32'h13020000;
          16'h0866 : blkif.rom_rdata <= 32'h97400000;
          16'h0867 : blkif.rom_rdata <= 32'h9380c002;
          16'h0868 : blkif.rom_rdata <= 32'h83a14000;
          16'h0869 : blkif.rom_rdata <= 32'h13830100;
          16'h086a : blkif.rom_rdata <= 32'hb71ef00f;
          16'h086b : blkif.rom_rdata <= 32'h938e0eff;
          16'h086c : blkif.rom_rdata <= 32'h6304d301;
          16'h086d : blkif.rom_rdata <= 32'h6f30805b;
          16'h086e : blkif.rom_rdata <= 32'h13021200;
          16'h086f : blkif.rom_rdata <= 32'h93022000;
          16'h0870 : blkif.rom_rdata <= 32'he31c52fc;
          16'h0871 : blkif.rom_rdata <= 32'h130ea014;
          16'h0872 : blkif.rom_rdata <= 32'h13020000;
          16'h0873 : blkif.rom_rdata <= 32'h97400000;
          16'h0874 : blkif.rom_rdata <= 32'h9380c0ff;
          16'h0875 : blkif.rom_rdata <= 32'h83a14000;
          16'h0876 : blkif.rom_rdata <= 32'h13000000;
          16'h0877 : blkif.rom_rdata <= 32'h13830100;
          16'h0878 : blkif.rom_rdata <= 32'hb7fe0ff0;
          16'h0879 : blkif.rom_rdata <= 32'h938efe00;
          16'h087a : blkif.rom_rdata <= 32'h6304d301;
          16'h087b : blkif.rom_rdata <= 32'h6f300058;
          16'h087c : blkif.rom_rdata <= 32'h13021200;
          16'h087d : blkif.rom_rdata <= 32'h93022000;
          16'h087e : blkif.rom_rdata <= 32'he31a52fc;
          16'h087f : blkif.rom_rdata <= 32'h130ec014;
          16'h0880 : blkif.rom_rdata <= 32'h13020000;
          16'h0881 : blkif.rom_rdata <= 32'h97400000;
          16'h0882 : blkif.rom_rdata <= 32'h938000fc;
          16'h0883 : blkif.rom_rdata <= 32'h83a14000;
          16'h0884 : blkif.rom_rdata <= 32'hb71ef00f;
          16'h0885 : blkif.rom_rdata <= 32'h938e0eff;
          16'h0886 : blkif.rom_rdata <= 32'h6384d101;
          16'h0887 : blkif.rom_rdata <= 32'h6f300055;
          16'h0888 : blkif.rom_rdata <= 32'h13021200;
          16'h0889 : blkif.rom_rdata <= 32'h93022000;
          16'h088a : blkif.rom_rdata <= 32'he31e52fc;
          16'h088b : blkif.rom_rdata <= 32'h130ee014;
          16'h088c : blkif.rom_rdata <= 32'h13020000;
          16'h088d : blkif.rom_rdata <= 32'h97400000;
          16'h088e : blkif.rom_rdata <= 32'h9380c0f8;
          16'h088f : blkif.rom_rdata <= 32'h13000000;
          16'h0890 : blkif.rom_rdata <= 32'h13000000;
          16'h0891 : blkif.rom_rdata <= 32'h83a14000;
          16'h0892 : blkif.rom_rdata <= 32'hb70e01ff;
          16'h0893 : blkif.rom_rdata <= 32'h938e0ef0;
          16'h0894 : blkif.rom_rdata <= 32'h6384d101;
          16'h0895 : blkif.rom_rdata <= 32'h6f308051;
          16'h0896 : blkif.rom_rdata <= 32'h13021200;
          16'h0897 : blkif.rom_rdata <= 32'h93022000;
          16'h0898 : blkif.rom_rdata <= 32'he31a52fc;
          16'h0899 : blkif.rom_rdata <= 32'hb7000080;
          16'h089a : blkif.rom_rdata <= 32'h93804000;
          16'h089b : blkif.rom_rdata <= 32'h1301f014;
          16'h089c : blkif.rom_rdata <= 32'h23a02000;
          16'h089d : blkif.rom_rdata <= 32'h97410000;
          16'h089e : blkif.rom_rdata <= 32'h9381c1f4;
          16'h089f : blkif.rom_rdata <= 32'h03a10100;
          16'h08a0 : blkif.rom_rdata <= 32'h13012000;
          16'h08a1 : blkif.rom_rdata <= 32'h930e2000;
          16'h08a2 : blkif.rom_rdata <= 32'h130ef014;
          16'h08a3 : blkif.rom_rdata <= 32'h6304d101;
          16'h08a4 : blkif.rom_rdata <= 32'h6f30c04d;
          16'h08a5 : blkif.rom_rdata <= 32'hb7000080;
          16'h08a6 : blkif.rom_rdata <= 32'h93804000;
          16'h08a7 : blkif.rom_rdata <= 32'h13010015;
          16'h08a8 : blkif.rom_rdata <= 32'h23a02000;
          16'h08a9 : blkif.rom_rdata <= 32'h97410000;
          16'h08aa : blkif.rom_rdata <= 32'h9381c1f1;
          16'h08ab : blkif.rom_rdata <= 32'h03a10100;
          16'h08ac : blkif.rom_rdata <= 32'h13000000;
          16'h08ad : blkif.rom_rdata <= 32'h13012000;
          16'h08ae : blkif.rom_rdata <= 32'h930e2000;
          16'h08af : blkif.rom_rdata <= 32'h130e0015;
          16'h08b0 : blkif.rom_rdata <= 32'h6304d101;
          16'h08b1 : blkif.rom_rdata <= 32'h6f30804a;
          16'h08b2 : blkif.rom_rdata <= 32'hb7000080;
          16'h08b3 : blkif.rom_rdata <= 32'h93804000;
          16'h08b4 : blkif.rom_rdata <= 32'h13011015;
          16'h08b5 : blkif.rom_rdata <= 32'h23a02000;
          16'h08b6 : blkif.rom_rdata <= 32'hb70001ff;
          16'h08b7 : blkif.rom_rdata <= 32'h938000f0;
          16'h08b8 : blkif.rom_rdata <= 32'h37110f0f;
          16'h08b9 : blkif.rom_rdata <= 32'h1301f1f0;
          16'h08ba : blkif.rom_rdata <= 32'hb3e12000;
          16'h08bb : blkif.rom_rdata <= 32'hb70e10ff;
          16'h08bc : blkif.rom_rdata <= 32'h938efef0;
          16'h08bd : blkif.rom_rdata <= 32'h130e1015;
          16'h08be : blkif.rom_rdata <= 32'h6384d101;
          16'h08bf : blkif.rom_rdata <= 32'h6f300047;
          16'h08c0 : blkif.rom_rdata <= 32'hb7000080;
          16'h08c1 : blkif.rom_rdata <= 32'h93804000;
          16'h08c2 : blkif.rom_rdata <= 32'h13014015;
          16'h08c3 : blkif.rom_rdata <= 32'h23a02000;
          16'h08c4 : blkif.rom_rdata <= 32'hb7f00ff0;
          16'h08c5 : blkif.rom_rdata <= 32'h9380f000;
          16'h08c6 : blkif.rom_rdata <= 32'h37f1f0f0;
          16'h08c7 : blkif.rom_rdata <= 32'h1301010f;
          16'h08c8 : blkif.rom_rdata <= 32'hb3e12000;
          16'h08c9 : blkif.rom_rdata <= 32'hb7fefff0;
          16'h08ca : blkif.rom_rdata <= 32'h938efe0f;
          16'h08cb : blkif.rom_rdata <= 32'h130e4015;
          16'h08cc : blkif.rom_rdata <= 32'h6384d101;
          16'h08cd : blkif.rom_rdata <= 32'h6f308043;
          16'h08ce : blkif.rom_rdata <= 32'hb7000080;
          16'h08cf : blkif.rom_rdata <= 32'h93804000;
          16'h08d0 : blkif.rom_rdata <= 32'h13015015;
          16'h08d1 : blkif.rom_rdata <= 32'h23a02000;
          16'h08d2 : blkif.rom_rdata <= 32'hb70001ff;
          16'h08d3 : blkif.rom_rdata <= 32'h938000f0;
          16'h08d4 : blkif.rom_rdata <= 32'h37110f0f;
          16'h08d5 : blkif.rom_rdata <= 32'h1301f1f0;
          16'h08d6 : blkif.rom_rdata <= 32'hb3e02000;
          16'h08d7 : blkif.rom_rdata <= 32'hb70e10ff;
          16'h08d8 : blkif.rom_rdata <= 32'h938efef0;
          16'h08d9 : blkif.rom_rdata <= 32'h130e5015;
          16'h08da : blkif.rom_rdata <= 32'h6384d001;
          16'h08db : blkif.rom_rdata <= 32'h6f300040;
          16'h08dc : blkif.rom_rdata <= 32'hb7000080;
          16'h08dd : blkif.rom_rdata <= 32'h93804000;
          16'h08de : blkif.rom_rdata <= 32'h13017015;
          16'h08df : blkif.rom_rdata <= 32'h23a02000;
          16'h08e0 : blkif.rom_rdata <= 32'hb70001ff;
          16'h08e1 : blkif.rom_rdata <= 32'h938000f0;
          16'h08e2 : blkif.rom_rdata <= 32'hb3e01000;
          16'h08e3 : blkif.rom_rdata <= 32'hb70e01ff;
          16'h08e4 : blkif.rom_rdata <= 32'h938e0ef0;
          16'h08e5 : blkif.rom_rdata <= 32'h130e7015;
          16'h08e6 : blkif.rom_rdata <= 32'h6384d001;
          16'h08e7 : blkif.rom_rdata <= 32'h6f30003d;
          16'h08e8 : blkif.rom_rdata <= 32'hb7000080;
          16'h08e9 : blkif.rom_rdata <= 32'h93804000;
          16'h08ea : blkif.rom_rdata <= 32'h13018015;
          16'h08eb : blkif.rom_rdata <= 32'h23a02000;
          16'h08ec : blkif.rom_rdata <= 32'h13020000;
          16'h08ed : blkif.rom_rdata <= 32'hb70001ff;
          16'h08ee : blkif.rom_rdata <= 32'h938000f0;
          16'h08ef : blkif.rom_rdata <= 32'h37110f0f;
          16'h08f0 : blkif.rom_rdata <= 32'h1301f1f0;
          16'h08f1 : blkif.rom_rdata <= 32'hb3e12000;
          16'h08f2 : blkif.rom_rdata <= 32'h13830100;
          16'h08f3 : blkif.rom_rdata <= 32'h13021200;
          16'h08f4 : blkif.rom_rdata <= 32'h93022000;
          16'h08f5 : blkif.rom_rdata <= 32'he31052fe;
          16'h08f6 : blkif.rom_rdata <= 32'hb70e10ff;
          16'h08f7 : blkif.rom_rdata <= 32'h938efef0;
          16'h08f8 : blkif.rom_rdata <= 32'h130e8015;
          16'h08f9 : blkif.rom_rdata <= 32'h6304d301;
          16'h08fa : blkif.rom_rdata <= 32'h6f304038;
          16'h08fb : blkif.rom_rdata <= 32'hb7000080;
          16'h08fc : blkif.rom_rdata <= 32'h93804000;
          16'h08fd : blkif.rom_rdata <= 32'h1301a015;
          16'h08fe : blkif.rom_rdata <= 32'h23a02000;
          16'h08ff : blkif.rom_rdata <= 32'h13020000;
          16'h0900 : blkif.rom_rdata <= 32'hb700ff00;
          16'h0901 : blkif.rom_rdata <= 32'h9380f00f;
          16'h0902 : blkif.rom_rdata <= 32'h37110f0f;
          16'h0903 : blkif.rom_rdata <= 32'h1301f1f0;
          16'h0904 : blkif.rom_rdata <= 32'hb3e12000;
          16'h0905 : blkif.rom_rdata <= 32'h13000000;
          16'h0906 : blkif.rom_rdata <= 32'h13000000;
          16'h0907 : blkif.rom_rdata <= 32'h13830100;
          16'h0908 : blkif.rom_rdata <= 32'h13021200;
          16'h0909 : blkif.rom_rdata <= 32'h93022000;
          16'h090a : blkif.rom_rdata <= 32'he31c52fc;
          16'h090b : blkif.rom_rdata <= 32'hb71eff0f;
          16'h090c : blkif.rom_rdata <= 32'h938efeff;
          16'h090d : blkif.rom_rdata <= 32'h130ea015;
          16'h090e : blkif.rom_rdata <= 32'h6304d301;
          16'h090f : blkif.rom_rdata <= 32'h6f300033;
          16'h0910 : blkif.rom_rdata <= 32'hb7000080;
          16'h0911 : blkif.rom_rdata <= 32'h93804000;
          16'h0912 : blkif.rom_rdata <= 32'h1301b015;
          16'h0913 : blkif.rom_rdata <= 32'h23a02000;
          16'h0914 : blkif.rom_rdata <= 32'h13020000;
          16'h0915 : blkif.rom_rdata <= 32'hb70001ff;
          16'h0916 : blkif.rom_rdata <= 32'h938000f0;
          16'h0917 : blkif.rom_rdata <= 32'h37110f0f;
          16'h0918 : blkif.rom_rdata <= 32'h1301f1f0;
          16'h0919 : blkif.rom_rdata <= 32'hb3e12000;
          16'h091a : blkif.rom_rdata <= 32'h13021200;
          16'h091b : blkif.rom_rdata <= 32'h93022000;
          16'h091c : blkif.rom_rdata <= 32'he31252fe;
          16'h091d : blkif.rom_rdata <= 32'hb70e10ff;
          16'h091e : blkif.rom_rdata <= 32'h938efef0;
          16'h091f : blkif.rom_rdata <= 32'h130eb015;
          16'h0920 : blkif.rom_rdata <= 32'h6384d101;
          16'h0921 : blkif.rom_rdata <= 32'h6f30802e;
          16'h0922 : blkif.rom_rdata <= 32'hb7000080;
          16'h0923 : blkif.rom_rdata <= 32'h93804000;
          16'h0924 : blkif.rom_rdata <= 32'h13010016;
          16'h0925 : blkif.rom_rdata <= 32'h23a02000;
          16'h0926 : blkif.rom_rdata <= 32'h13020000;
          16'h0927 : blkif.rom_rdata <= 32'hb700ff00;
          16'h0928 : blkif.rom_rdata <= 32'h9380f00f;
          16'h0929 : blkif.rom_rdata <= 32'h13000000;
          16'h092a : blkif.rom_rdata <= 32'h13000000;
          16'h092b : blkif.rom_rdata <= 32'h37110f0f;
          16'h092c : blkif.rom_rdata <= 32'h1301f1f0;
          16'h092d : blkif.rom_rdata <= 32'hb3e12000;
          16'h092e : blkif.rom_rdata <= 32'h13021200;
          16'h092f : blkif.rom_rdata <= 32'h93022000;
          16'h0930 : blkif.rom_rdata <= 32'he31e52fc;
          16'h0931 : blkif.rom_rdata <= 32'hb71eff0f;
          16'h0932 : blkif.rom_rdata <= 32'h938efeff;
          16'h0933 : blkif.rom_rdata <= 32'h130e0016;
          16'h0934 : blkif.rom_rdata <= 32'h6384d101;
          16'h0935 : blkif.rom_rdata <= 32'h6f308029;
          16'h0936 : blkif.rom_rdata <= 32'hb7000080;
          16'h0937 : blkif.rom_rdata <= 32'h93804000;
          16'h0938 : blkif.rom_rdata <= 32'h13011016;
          16'h0939 : blkif.rom_rdata <= 32'h23a02000;
          16'h093a : blkif.rom_rdata <= 32'h13020000;
          16'h093b : blkif.rom_rdata <= 32'h37110f0f;
          16'h093c : blkif.rom_rdata <= 32'h1301f1f0;
          16'h093d : blkif.rom_rdata <= 32'hb70001ff;
          16'h093e : blkif.rom_rdata <= 32'h938000f0;
          16'h093f : blkif.rom_rdata <= 32'hb3e12000;
          16'h0940 : blkif.rom_rdata <= 32'h13021200;
          16'h0941 : blkif.rom_rdata <= 32'h93022000;
          16'h0942 : blkif.rom_rdata <= 32'he31252fe;
          16'h0943 : blkif.rom_rdata <= 32'hb70e10ff;
          16'h0944 : blkif.rom_rdata <= 32'h938efef0;
          16'h0945 : blkif.rom_rdata <= 32'h130e1016;
          16'h0946 : blkif.rom_rdata <= 32'h6384d101;
          16'h0947 : blkif.rom_rdata <= 32'h6f300025;
          16'h0948 : blkif.rom_rdata <= 32'hb7000080;
          16'h0949 : blkif.rom_rdata <= 32'h93804000;
          16'h094a : blkif.rom_rdata <= 32'h13016016;
          16'h094b : blkif.rom_rdata <= 32'h23a02000;
          16'h094c : blkif.rom_rdata <= 32'h13020000;
          16'h094d : blkif.rom_rdata <= 32'h37110f0f;
          16'h094e : blkif.rom_rdata <= 32'h1301f1f0;
          16'h094f : blkif.rom_rdata <= 32'h13000000;
          16'h0950 : blkif.rom_rdata <= 32'h13000000;
          16'h0951 : blkif.rom_rdata <= 32'hb700ff00;
          16'h0952 : blkif.rom_rdata <= 32'h9380f00f;
          16'h0953 : blkif.rom_rdata <= 32'hb3e12000;
          16'h0954 : blkif.rom_rdata <= 32'h13021200;
          16'h0955 : blkif.rom_rdata <= 32'h93022000;
          16'h0956 : blkif.rom_rdata <= 32'he31e52fc;
          16'h0957 : blkif.rom_rdata <= 32'hb71eff0f;
          16'h0958 : blkif.rom_rdata <= 32'h938efeff;
          16'h0959 : blkif.rom_rdata <= 32'h130e6016;
          16'h095a : blkif.rom_rdata <= 32'h6384d101;
          16'h095b : blkif.rom_rdata <= 32'h6f300020;
          16'h095c : blkif.rom_rdata <= 32'hb7000080;
          16'h095d : blkif.rom_rdata <= 32'h93804000;
          16'h095e : blkif.rom_rdata <= 32'h13017016;
          16'h095f : blkif.rom_rdata <= 32'h23a02000;
          16'h0960 : blkif.rom_rdata <= 32'hb70001ff;
          16'h0961 : blkif.rom_rdata <= 32'h938000f0;
          16'h0962 : blkif.rom_rdata <= 32'h33611000;
          16'h0963 : blkif.rom_rdata <= 32'hb70e01ff;
          16'h0964 : blkif.rom_rdata <= 32'h938e0ef0;
          16'h0965 : blkif.rom_rdata <= 32'h130e7016;
          16'h0966 : blkif.rom_rdata <= 32'h6304d101;
          16'h0967 : blkif.rom_rdata <= 32'h6f30001d;
          16'h0968 : blkif.rom_rdata <= 32'hb7000080;
          16'h0969 : blkif.rom_rdata <= 32'h93804000;
          16'h096a : blkif.rom_rdata <= 32'h13019016;
          16'h096b : blkif.rom_rdata <= 32'h23a02000;
          16'h096c : blkif.rom_rdata <= 32'hb3600000;
          16'h096d : blkif.rom_rdata <= 32'h930e0000;
          16'h096e : blkif.rom_rdata <= 32'h130e9016;
          16'h096f : blkif.rom_rdata <= 32'h6384d001;
          16'h0970 : blkif.rom_rdata <= 32'h6f30c01a;
          16'h0971 : blkif.rom_rdata <= 32'hb7000080;
          16'h0972 : blkif.rom_rdata <= 32'h93804000;
          16'h0973 : blkif.rom_rdata <= 32'h1301a016;
          16'h0974 : blkif.rom_rdata <= 32'h23a02000;
          16'h0975 : blkif.rom_rdata <= 32'hb7101111;
          16'h0976 : blkif.rom_rdata <= 32'h93801011;
          16'h0977 : blkif.rom_rdata <= 32'h37212222;
          16'h0978 : blkif.rom_rdata <= 32'h13012122;
          16'h0979 : blkif.rom_rdata <= 32'h33e02000;
          16'h097a : blkif.rom_rdata <= 32'h930e0000;
          16'h097b : blkif.rom_rdata <= 32'h130ea016;
          16'h097c : blkif.rom_rdata <= 32'h6304d001;
          16'h097d : blkif.rom_rdata <= 32'h6f308017;
          16'h097e : blkif.rom_rdata <= 32'hb7000080;
          16'h097f : blkif.rom_rdata <= 32'h93804000;
          16'h0980 : blkif.rom_rdata <= 32'h1301b016;
          16'h0981 : blkif.rom_rdata <= 32'h23a02000;
          16'h0982 : blkif.rom_rdata <= 32'hb70001ff;
          16'h0983 : blkif.rom_rdata <= 32'h938000f0;
          16'h0984 : blkif.rom_rdata <= 32'h93e1f0f0;
          16'h0985 : blkif.rom_rdata <= 32'h930ef0f0;
          16'h0986 : blkif.rom_rdata <= 32'h130eb016;
          16'h0987 : blkif.rom_rdata <= 32'h6384d101;
          16'h0988 : blkif.rom_rdata <= 32'h6f30c014;
          16'h0989 : blkif.rom_rdata <= 32'hb7000080;
          16'h098a : blkif.rom_rdata <= 32'h93804000;
          16'h098b : blkif.rom_rdata <= 32'h1301e016;
          16'h098c : blkif.rom_rdata <= 32'h23a02000;
          16'h098d : blkif.rom_rdata <= 32'hb7f00ff0;
          16'h098e : blkif.rom_rdata <= 32'h9380f000;
          16'h098f : blkif.rom_rdata <= 32'h93e1000f;
          16'h0990 : blkif.rom_rdata <= 32'hb7fe0ff0;
          16'h0991 : blkif.rom_rdata <= 32'h938efe0f;
          16'h0992 : blkif.rom_rdata <= 32'h130ee016;
          16'h0993 : blkif.rom_rdata <= 32'h6384d101;
          16'h0994 : blkif.rom_rdata <= 32'h6f30c011;
          16'h0995 : blkif.rom_rdata <= 32'hb7000080;
          16'h0996 : blkif.rom_rdata <= 32'h93804000;
          16'h0997 : blkif.rom_rdata <= 32'h1301f016;
          16'h0998 : blkif.rom_rdata <= 32'h23a02000;
          16'h0999 : blkif.rom_rdata <= 32'hb70001ff;
          16'h099a : blkif.rom_rdata <= 32'h938000f0;
          16'h099b : blkif.rom_rdata <= 32'h93e0000f;
          16'h099c : blkif.rom_rdata <= 32'hb70e01ff;
          16'h099d : blkif.rom_rdata <= 32'h938e0eff;
          16'h099e : blkif.rom_rdata <= 32'h130ef016;
          16'h099f : blkif.rom_rdata <= 32'h6384d001;
          16'h09a0 : blkif.rom_rdata <= 32'h6f30c00e;
          16'h09a1 : blkif.rom_rdata <= 32'hb7000080;
          16'h09a2 : blkif.rom_rdata <= 32'h93804000;
          16'h09a3 : blkif.rom_rdata <= 32'h13011017;
          16'h09a4 : blkif.rom_rdata <= 32'h23a02000;
          16'h09a5 : blkif.rom_rdata <= 32'h13020000;
          16'h09a6 : blkif.rom_rdata <= 32'hb700ff00;
          16'h09a7 : blkif.rom_rdata <= 32'h9380f00f;
          16'h09a8 : blkif.rom_rdata <= 32'h93e1f070;
          16'h09a9 : blkif.rom_rdata <= 32'h13000000;
          16'h09aa : blkif.rom_rdata <= 32'h13830100;
          16'h09ab : blkif.rom_rdata <= 32'h13021200;
          16'h09ac : blkif.rom_rdata <= 32'h93022000;
          16'h09ad : blkif.rom_rdata <= 32'he31252fe;
          16'h09ae : blkif.rom_rdata <= 32'hb70eff00;
          16'h09af : blkif.rom_rdata <= 32'h938efe7f;
          16'h09b0 : blkif.rom_rdata <= 32'h130e1017;
          16'h09b1 : blkif.rom_rdata <= 32'h6304d301;
          16'h09b2 : blkif.rom_rdata <= 32'h6f30400a;
          16'h09b3 : blkif.rom_rdata <= 32'hb7000080;
          16'h09b4 : blkif.rom_rdata <= 32'h93804000;
          16'h09b5 : blkif.rom_rdata <= 32'h13012017;
          16'h09b6 : blkif.rom_rdata <= 32'h23a02000;
          16'h09b7 : blkif.rom_rdata <= 32'h13020000;
          16'h09b8 : blkif.rom_rdata <= 32'hb7f00ff0;
          16'h09b9 : blkif.rom_rdata <= 32'h9380f000;
          16'h09ba : blkif.rom_rdata <= 32'h93e1000f;
          16'h09bb : blkif.rom_rdata <= 32'h13000000;
          16'h09bc : blkif.rom_rdata <= 32'h13000000;
          16'h09bd : blkif.rom_rdata <= 32'h13830100;
          16'h09be : blkif.rom_rdata <= 32'h13021200;
          16'h09bf : blkif.rom_rdata <= 32'h93022000;
          16'h09c0 : blkif.rom_rdata <= 32'he31052fe;
          16'h09c1 : blkif.rom_rdata <= 32'hb7fe0ff0;
          16'h09c2 : blkif.rom_rdata <= 32'h938efe0f;
          16'h09c3 : blkif.rom_rdata <= 32'h130e2017;
          16'h09c4 : blkif.rom_rdata <= 32'h6304d301;
          16'h09c5 : blkif.rom_rdata <= 32'h6f308005;
          16'h09c6 : blkif.rom_rdata <= 32'hb7000080;
          16'h09c7 : blkif.rom_rdata <= 32'h93804000;
          16'h09c8 : blkif.rom_rdata <= 32'h13013017;
          16'h09c9 : blkif.rom_rdata <= 32'h23a02000;
          16'h09ca : blkif.rom_rdata <= 32'h13020000;
          16'h09cb : blkif.rom_rdata <= 32'hb710f00f;
          16'h09cc : blkif.rom_rdata <= 32'h938000ff;
          16'h09cd : blkif.rom_rdata <= 32'h93e1000f;
          16'h09ce : blkif.rom_rdata <= 32'h13021200;
          16'h09cf : blkif.rom_rdata <= 32'h93022000;
          16'h09d0 : blkif.rom_rdata <= 32'he31652fe;
          16'h09d1 : blkif.rom_rdata <= 32'hb71ef00f;
          16'h09d2 : blkif.rom_rdata <= 32'h938e0eff;
          16'h09d3 : blkif.rom_rdata <= 32'h130e3017;
          16'h09d4 : blkif.rom_rdata <= 32'h6384d101;
          16'h09d5 : blkif.rom_rdata <= 32'h6f308001;
          16'h09d6 : blkif.rom_rdata <= 32'hb7000080;
          16'h09d7 : blkif.rom_rdata <= 32'h93804000;
          16'h09d8 : blkif.rom_rdata <= 32'h13015017;
          16'h09d9 : blkif.rom_rdata <= 32'h23a02000;
          16'h09da : blkif.rom_rdata <= 32'h13020000;
          16'h09db : blkif.rom_rdata <= 32'hb7f00ff0;
          16'h09dc : blkif.rom_rdata <= 32'h9380f000;
          16'h09dd : blkif.rom_rdata <= 32'h13000000;
          16'h09de : blkif.rom_rdata <= 32'h13000000;
          16'h09df : blkif.rom_rdata <= 32'h93e1000f;
          16'h09e0 : blkif.rom_rdata <= 32'h13021200;
          16'h09e1 : blkif.rom_rdata <= 32'h93022000;
          16'h09e2 : blkif.rom_rdata <= 32'he31252fe;
          16'h09e3 : blkif.rom_rdata <= 32'hb7fe0ff0;
          16'h09e4 : blkif.rom_rdata <= 32'h938efe0f;
          16'h09e5 : blkif.rom_rdata <= 32'h130e5017;
          16'h09e6 : blkif.rom_rdata <= 32'h6384d101;
          16'h09e7 : blkif.rom_rdata <= 32'h6f20107d;
          16'h09e8 : blkif.rom_rdata <= 32'hb7000080;
          16'h09e9 : blkif.rom_rdata <= 32'h93804000;
          16'h09ea : blkif.rom_rdata <= 32'h13016017;
          16'h09eb : blkif.rom_rdata <= 32'h23a02000;
          16'h09ec : blkif.rom_rdata <= 32'h9360000f;
          16'h09ed : blkif.rom_rdata <= 32'h930e000f;
          16'h09ee : blkif.rom_rdata <= 32'h130e6017;
          16'h09ef : blkif.rom_rdata <= 32'h6384d001;
          16'h09f0 : blkif.rom_rdata <= 32'h6f20d07a;
          16'h09f1 : blkif.rom_rdata <= 32'hb7000080;
          16'h09f2 : blkif.rom_rdata <= 32'h93804000;
          16'h09f3 : blkif.rom_rdata <= 32'h13017017;
          16'h09f4 : blkif.rom_rdata <= 32'h23a02000;
          16'h09f5 : blkif.rom_rdata <= 32'hb700ff00;
          16'h09f6 : blkif.rom_rdata <= 32'h9380f00f;
          16'h09f7 : blkif.rom_rdata <= 32'h13e0f070;
          16'h09f8 : blkif.rom_rdata <= 32'h930e0000;
          16'h09f9 : blkif.rom_rdata <= 32'h130e7017;
          16'h09fa : blkif.rom_rdata <= 32'h6304d001;
          16'h09fb : blkif.rom_rdata <= 32'h6f201078;
          16'h09fc : blkif.rom_rdata <= 32'hb7f0efef;
          16'h09fd : blkif.rom_rdata <= 32'h9380f0fe;
          16'h09fe : blkif.rom_rdata <= 32'h17610000;
          16'h09ff : blkif.rom_rdata <= 32'h13018180;
          16'h0a00 : blkif.rom_rdata <= 32'h23201100;
          16'h0a01 : blkif.rom_rdata <= 32'h23221100;
          16'h0a02 : blkif.rom_rdata <= 32'h23241100;
          16'h0a03 : blkif.rom_rdata <= 32'hb7000080;
          16'h0a04 : blkif.rom_rdata <= 32'h93804000;
          16'h0a05 : blkif.rom_rdata <= 32'h13018017;
          16'h0a06 : blkif.rom_rdata <= 32'h23a02000;
          16'h0a07 : blkif.rom_rdata <= 32'h97500000;
          16'h0a08 : blkif.rom_rdata <= 32'h9380407e;
          16'h0a09 : blkif.rom_rdata <= 32'h1301a0fa;
          16'h0a0a : blkif.rom_rdata <= 32'h23802000;
          16'h0a0b : blkif.rom_rdata <= 32'h83810000;
          16'h0a0c : blkif.rom_rdata <= 32'h930ea0fa;
          16'h0a0d : blkif.rom_rdata <= 32'h130e8017;
          16'h0a0e : blkif.rom_rdata <= 32'h6384d101;
          16'h0a0f : blkif.rom_rdata <= 32'h6f201073;
          16'h0a10 : blkif.rom_rdata <= 32'hb7000080;
          16'h0a11 : blkif.rom_rdata <= 32'h93804000;
          16'h0a12 : blkif.rom_rdata <= 32'h13019017;
          16'h0a13 : blkif.rom_rdata <= 32'h23a02000;
          16'h0a14 : blkif.rom_rdata <= 32'h97500000;
          16'h0a15 : blkif.rom_rdata <= 32'h9380007b;
          16'h0a16 : blkif.rom_rdata <= 32'h13010000;
          16'h0a17 : blkif.rom_rdata <= 32'ha3802000;
          16'h0a18 : blkif.rom_rdata <= 32'h83811000;
          16'h0a19 : blkif.rom_rdata <= 32'h930e0000;
          16'h0a1a : blkif.rom_rdata <= 32'h130e9017;
          16'h0a1b : blkif.rom_rdata <= 32'h6384d101;
          16'h0a1c : blkif.rom_rdata <= 32'h6f20d06f;
          16'h0a1d : blkif.rom_rdata <= 32'hb7000080;
          16'h0a1e : blkif.rom_rdata <= 32'h93804000;
          16'h0a1f : blkif.rom_rdata <= 32'h1301a017;
          16'h0a20 : blkif.rom_rdata <= 32'h23a02000;
          16'h0a21 : blkif.rom_rdata <= 32'h97500000;
          16'h0a22 : blkif.rom_rdata <= 32'h9380c077;
          16'h0a23 : blkif.rom_rdata <= 32'h37f1ffff;
          16'h0a24 : blkif.rom_rdata <= 32'h130101fa;
          16'h0a25 : blkif.rom_rdata <= 32'h23812000;
          16'h0a26 : blkif.rom_rdata <= 32'h83912000;
          16'h0a27 : blkif.rom_rdata <= 32'hb7feffff;
          16'h0a28 : blkif.rom_rdata <= 32'h938e0efa;
          16'h0a29 : blkif.rom_rdata <= 32'h130ea017;
          16'h0a2a : blkif.rom_rdata <= 32'h6384d101;
          16'h0a2b : blkif.rom_rdata <= 32'h6f20106c;
          16'h0a2c : blkif.rom_rdata <= 32'hb7000080;
          16'h0a2d : blkif.rom_rdata <= 32'h93804000;
          16'h0a2e : blkif.rom_rdata <= 32'h1301c017;
          16'h0a2f : blkif.rom_rdata <= 32'h23a02000;
          16'h0a30 : blkif.rom_rdata <= 32'h97500000;
          16'h0a31 : blkif.rom_rdata <= 32'h93800074;
          16'h0a32 : blkif.rom_rdata <= 32'h1301a000;
          16'h0a33 : blkif.rom_rdata <= 32'ha3812000;
          16'h0a34 : blkif.rom_rdata <= 32'h83813000;
          16'h0a35 : blkif.rom_rdata <= 32'h930ea000;
          16'h0a36 : blkif.rom_rdata <= 32'h130ec017;
          16'h0a37 : blkif.rom_rdata <= 32'h6384d101;
          16'h0a38 : blkif.rom_rdata <= 32'h6f20d068;
          16'h0a39 : blkif.rom_rdata <= 32'hb7000080;
          16'h0a3a : blkif.rom_rdata <= 32'h93804000;
          16'h0a3b : blkif.rom_rdata <= 32'h1301d017;
          16'h0a3c : blkif.rom_rdata <= 32'h23a02000;
          16'h0a3d : blkif.rom_rdata <= 32'h97500000;
          16'h0a3e : blkif.rom_rdata <= 32'h93803071;
          16'h0a3f : blkif.rom_rdata <= 32'h1301a0fa;
          16'h0a40 : blkif.rom_rdata <= 32'ha38e20fe;
          16'h0a41 : blkif.rom_rdata <= 32'h8381d0ff;
          16'h0a42 : blkif.rom_rdata <= 32'h930ea0fa;
          16'h0a43 : blkif.rom_rdata <= 32'h130ed017;
          16'h0a44 : blkif.rom_rdata <= 32'h6384d101;
          16'h0a45 : blkif.rom_rdata <= 32'h6f209065;
          16'h0a46 : blkif.rom_rdata <= 32'hb7000080;
          16'h0a47 : blkif.rom_rdata <= 32'h93804000;
          16'h0a48 : blkif.rom_rdata <= 32'h1301e017;
          16'h0a49 : blkif.rom_rdata <= 32'h23a02000;
          16'h0a4a : blkif.rom_rdata <= 32'h97500000;
          16'h0a4b : blkif.rom_rdata <= 32'h9380f06d;
          16'h0a4c : blkif.rom_rdata <= 32'h13010000;
          16'h0a4d : blkif.rom_rdata <= 32'h238f20fe;
          16'h0a4e : blkif.rom_rdata <= 32'h8381e0ff;
          16'h0a4f : blkif.rom_rdata <= 32'h930e0000;
          16'h0a50 : blkif.rom_rdata <= 32'h130ee017;
          16'h0a51 : blkif.rom_rdata <= 32'h6384d101;
          16'h0a52 : blkif.rom_rdata <= 32'h6f205062;
          16'h0a53 : blkif.rom_rdata <= 32'hb7000080;
          16'h0a54 : blkif.rom_rdata <= 32'h93804000;
          16'h0a55 : blkif.rom_rdata <= 32'h13010018;
          16'h0a56 : blkif.rom_rdata <= 32'h23a02000;
          16'h0a57 : blkif.rom_rdata <= 32'h97500000;
          16'h0a58 : blkif.rom_rdata <= 32'h9380b06a;
          16'h0a59 : blkif.rom_rdata <= 32'h1301a000;
          16'h0a5a : blkif.rom_rdata <= 32'h23802000;
          16'h0a5b : blkif.rom_rdata <= 32'h83810000;
          16'h0a5c : blkif.rom_rdata <= 32'h930ea000;
          16'h0a5d : blkif.rom_rdata <= 32'h130e0018;
          16'h0a5e : blkif.rom_rdata <= 32'h6384d101;
          16'h0a5f : blkif.rom_rdata <= 32'h6f20105f;
          16'h0a60 : blkif.rom_rdata <= 32'hb7000080;
          16'h0a61 : blkif.rom_rdata <= 32'h93804000;
          16'h0a62 : blkif.rom_rdata <= 32'h13011018;
          16'h0a63 : blkif.rom_rdata <= 32'h23a02000;
          16'h0a64 : blkif.rom_rdata <= 32'h97500000;
          16'h0a65 : blkif.rom_rdata <= 32'h93808067;
          16'h0a66 : blkif.rom_rdata <= 32'h37513412;
          16'h0a67 : blkif.rom_rdata <= 32'h13018167;
          16'h0a68 : blkif.rom_rdata <= 32'h138200fe;
          16'h0a69 : blkif.rom_rdata <= 32'h23002202;
          16'h0a6a : blkif.rom_rdata <= 32'h83810000;
          16'h0a6b : blkif.rom_rdata <= 32'h930e8007;
          16'h0a6c : blkif.rom_rdata <= 32'h130e1018;
          16'h0a6d : blkif.rom_rdata <= 32'h6384d101;
          16'h0a6e : blkif.rom_rdata <= 32'h6f20505b;
          16'h0a6f : blkif.rom_rdata <= 32'hb7000080;
          16'h0a70 : blkif.rom_rdata <= 32'h93804000;
          16'h0a71 : blkif.rom_rdata <= 32'h13012018;
          16'h0a72 : blkif.rom_rdata <= 32'h23a02000;
          16'h0a73 : blkif.rom_rdata <= 32'h97500000;
          16'h0a74 : blkif.rom_rdata <= 32'h9380c063;
          16'h0a75 : blkif.rom_rdata <= 32'h37310000;
          16'h0a76 : blkif.rom_rdata <= 32'h13018109;
          16'h0a77 : blkif.rom_rdata <= 32'h9380a0ff;
          16'h0a78 : blkif.rom_rdata <= 32'ha3832000;
          16'h0a79 : blkif.rom_rdata <= 32'h17520000;
          16'h0a7a : blkif.rom_rdata <= 32'h13025262;
          16'h0a7b : blkif.rom_rdata <= 32'h83010200;
          16'h0a7c : blkif.rom_rdata <= 32'h930e80f9;
          16'h0a7d : blkif.rom_rdata <= 32'h130e2018;
          16'h0a7e : blkif.rom_rdata <= 32'h6384d101;
          16'h0a7f : blkif.rom_rdata <= 32'h6f201057;
          16'h0a80 : blkif.rom_rdata <= 32'h130e3018;
          16'h0a81 : blkif.rom_rdata <= 32'h13020000;
          16'h0a82 : blkif.rom_rdata <= 32'h9300d0fd;
          16'h0a83 : blkif.rom_rdata <= 32'h17510000;
          16'h0a84 : blkif.rom_rdata <= 32'h1301415f;
          16'h0a85 : blkif.rom_rdata <= 32'h23001100;
          16'h0a86 : blkif.rom_rdata <= 32'h83010100;
          16'h0a87 : blkif.rom_rdata <= 32'h930ed0fd;
          16'h0a88 : blkif.rom_rdata <= 32'h6384d101;
          16'h0a89 : blkif.rom_rdata <= 32'h6f209054;
          16'h0a8a : blkif.rom_rdata <= 32'h13021200;
          16'h0a8b : blkif.rom_rdata <= 32'h93022000;
          16'h0a8c : blkif.rom_rdata <= 32'he31c52fc;
          16'h0a8d : blkif.rom_rdata <= 32'h130e4018;
          16'h0a8e : blkif.rom_rdata <= 32'h13020000;
          16'h0a8f : blkif.rom_rdata <= 32'h9300d0fc;
          16'h0a90 : blkif.rom_rdata <= 32'h17510000;
          16'h0a91 : blkif.rom_rdata <= 32'h1301015c;
          16'h0a92 : blkif.rom_rdata <= 32'h13000000;
          16'h0a93 : blkif.rom_rdata <= 32'ha3001100;
          16'h0a94 : blkif.rom_rdata <= 32'h83011100;
          16'h0a95 : blkif.rom_rdata <= 32'h930ed0fc;
          16'h0a96 : blkif.rom_rdata <= 32'h6384d101;
          16'h0a97 : blkif.rom_rdata <= 32'h6f201051;
          16'h0a98 : blkif.rom_rdata <= 32'h13021200;
          16'h0a99 : blkif.rom_rdata <= 32'h93022000;
          16'h0a9a : blkif.rom_rdata <= 32'he31a52fc;
          16'h0a9b : blkif.rom_rdata <= 32'h130e7018;
          16'h0a9c : blkif.rom_rdata <= 32'h13020000;
          16'h0a9d : blkif.rom_rdata <= 32'h9300b0fb;
          16'h0a9e : blkif.rom_rdata <= 32'h13000000;
          16'h0a9f : blkif.rom_rdata <= 32'h17510000;
          16'h0aa0 : blkif.rom_rdata <= 32'h13014158;
          16'h0aa1 : blkif.rom_rdata <= 32'h13000000;
          16'h0aa2 : blkif.rom_rdata <= 32'h23021100;
          16'h0aa3 : blkif.rom_rdata <= 32'h83014100;
          16'h0aa4 : blkif.rom_rdata <= 32'h930eb0fb;
          16'h0aa5 : blkif.rom_rdata <= 32'h6384d101;
          16'h0aa6 : blkif.rom_rdata <= 32'h6f20504d;
          16'h0aa7 : blkif.rom_rdata <= 32'h13021200;
          16'h0aa8 : blkif.rom_rdata <= 32'h93022000;
          16'h0aa9 : blkif.rom_rdata <= 32'he31852fc;
          16'h0aaa : blkif.rom_rdata <= 32'h130e9018;
          16'h0aab : blkif.rom_rdata <= 32'h13020000;
          16'h0aac : blkif.rom_rdata <= 32'h17510000;
          16'h0aad : blkif.rom_rdata <= 32'h13010155;
          16'h0aae : blkif.rom_rdata <= 32'h93003003;
          16'h0aaf : blkif.rom_rdata <= 32'h23001100;
          16'h0ab0 : blkif.rom_rdata <= 32'h83010100;
          16'h0ab1 : blkif.rom_rdata <= 32'h930e3003;
          16'h0ab2 : blkif.rom_rdata <= 32'h6384d101;
          16'h0ab3 : blkif.rom_rdata <= 32'h6f20104a;
          16'h0ab4 : blkif.rom_rdata <= 32'h13021200;
          16'h0ab5 : blkif.rom_rdata <= 32'h93022000;
          16'h0ab6 : blkif.rom_rdata <= 32'he31c52fc;
          16'h0ab7 : blkif.rom_rdata <= 32'h130ea018;
          16'h0ab8 : blkif.rom_rdata <= 32'h13020000;
          16'h0ab9 : blkif.rom_rdata <= 32'h17510000;
          16'h0aba : blkif.rom_rdata <= 32'h1301c151;
          16'h0abb : blkif.rom_rdata <= 32'h93003002;
          16'h0abc : blkif.rom_rdata <= 32'h13000000;
          16'h0abd : blkif.rom_rdata <= 32'ha3001100;
          16'h0abe : blkif.rom_rdata <= 32'h83011100;
          16'h0abf : blkif.rom_rdata <= 32'h930e3002;
          16'h0ac0 : blkif.rom_rdata <= 32'h6384d101;
          16'h0ac1 : blkif.rom_rdata <= 32'h6f209046;
          16'h0ac2 : blkif.rom_rdata <= 32'h13021200;
          16'h0ac3 : blkif.rom_rdata <= 32'h93022000;
          16'h0ac4 : blkif.rom_rdata <= 32'he31a52fc;
          16'h0ac5 : blkif.rom_rdata <= 32'h1305f00e;
          16'h0ac6 : blkif.rom_rdata <= 32'h97550000;
          16'h0ac7 : blkif.rom_rdata <= 32'h9385854e;
          16'h0ac8 : blkif.rom_rdata <= 32'ha381a500;
          16'h0ac9 : blkif.rom_rdata <= 32'hb7c0efbe;
          16'h0aca : blkif.rom_rdata <= 32'h9380f0ee;
          16'h0acb : blkif.rom_rdata <= 32'h17510000;
          16'h0acc : blkif.rom_rdata <= 32'h1301414e;
          16'h0acd : blkif.rom_rdata <= 32'h23201100;
          16'h0ace : blkif.rom_rdata <= 32'h23221100;
          16'h0acf : blkif.rom_rdata <= 32'h23241100;
          16'h0ad0 : blkif.rom_rdata <= 32'h23261100;
          16'h0ad1 : blkif.rom_rdata <= 32'h23281100;
          16'h0ad2 : blkif.rom_rdata <= 32'hb7000080;
          16'h0ad3 : blkif.rom_rdata <= 32'h93804000;
          16'h0ad4 : blkif.rom_rdata <= 32'h1301f018;
          16'h0ad5 : blkif.rom_rdata <= 32'h23a02000;
          16'h0ad6 : blkif.rom_rdata <= 32'h97500000;
          16'h0ad7 : blkif.rom_rdata <= 32'h9380804b;
          16'h0ad8 : blkif.rom_rdata <= 32'h1301a00a;
          16'h0ad9 : blkif.rom_rdata <= 32'h23902000;
          16'h0ada : blkif.rom_rdata <= 32'h83910000;
          16'h0adb : blkif.rom_rdata <= 32'h930ea00a;
          16'h0adc : blkif.rom_rdata <= 32'h130ef018;
          16'h0add : blkif.rom_rdata <= 32'h6384d101;
          16'h0ade : blkif.rom_rdata <= 32'h6f20503f;
          16'h0adf : blkif.rom_rdata <= 32'hb7000080;
          16'h0ae0 : blkif.rom_rdata <= 32'h93804000;
          16'h0ae1 : blkif.rom_rdata <= 32'h13010019;
          16'h0ae2 : blkif.rom_rdata <= 32'h23a02000;
          16'h0ae3 : blkif.rom_rdata <= 32'h97500000;
          16'h0ae4 : blkif.rom_rdata <= 32'h93804048;
          16'h0ae5 : blkif.rom_rdata <= 32'h37b1ffff;
          16'h0ae6 : blkif.rom_rdata <= 32'h130101a0;
          16'h0ae7 : blkif.rom_rdata <= 32'h23912000;
          16'h0ae8 : blkif.rom_rdata <= 32'h83912000;
          16'h0ae9 : blkif.rom_rdata <= 32'hb7beffff;
          16'h0aea : blkif.rom_rdata <= 32'h938e0ea0;
          16'h0aeb : blkif.rom_rdata <= 32'h130e0019;
          16'h0aec : blkif.rom_rdata <= 32'h6384d101;
          16'h0aed : blkif.rom_rdata <= 32'h6f20903b;
          16'h0aee : blkif.rom_rdata <= 32'hb7000080;
          16'h0aef : blkif.rom_rdata <= 32'h93804000;
          16'h0af0 : blkif.rom_rdata <= 32'h13011019;
          16'h0af1 : blkif.rom_rdata <= 32'h23a02000;
          16'h0af2 : blkif.rom_rdata <= 32'h97500000;
          16'h0af3 : blkif.rom_rdata <= 32'h93808044;
          16'h0af4 : blkif.rom_rdata <= 32'h3711efbe;
          16'h0af5 : blkif.rom_rdata <= 32'h130101aa;
          16'h0af6 : blkif.rom_rdata <= 32'h23922000;
          16'h0af7 : blkif.rom_rdata <= 32'h83a14000;
          16'h0af8 : blkif.rom_rdata <= 32'hb71eefbe;
          16'h0af9 : blkif.rom_rdata <= 32'h938e0eaa;
          16'h0afa : blkif.rom_rdata <= 32'h130e1019;
          16'h0afb : blkif.rom_rdata <= 32'h6384d101;
          16'h0afc : blkif.rom_rdata <= 32'h6f20d037;
          16'h0afd : blkif.rom_rdata <= 32'hb7000080;
          16'h0afe : blkif.rom_rdata <= 32'h93804000;
          16'h0aff : blkif.rom_rdata <= 32'h13012019;
          16'h0b00 : blkif.rom_rdata <= 32'h23a02000;
          16'h0b01 : blkif.rom_rdata <= 32'h97500000;
          16'h0b02 : blkif.rom_rdata <= 32'h9380c040;
          16'h0b03 : blkif.rom_rdata <= 32'h37a1ffff;
          16'h0b04 : blkif.rom_rdata <= 32'h1301a100;
          16'h0b05 : blkif.rom_rdata <= 32'h23932000;
          16'h0b06 : blkif.rom_rdata <= 32'h83916000;
          16'h0b07 : blkif.rom_rdata <= 32'hb7aeffff;
          16'h0b08 : blkif.rom_rdata <= 32'h938eae00;
          16'h0b09 : blkif.rom_rdata <= 32'h130e2019;
          16'h0b0a : blkif.rom_rdata <= 32'h6384d101;
          16'h0b0b : blkif.rom_rdata <= 32'h6f201034;
          16'h0b0c : blkif.rom_rdata <= 32'hb7000080;
          16'h0b0d : blkif.rom_rdata <= 32'h93804000;
          16'h0b0e : blkif.rom_rdata <= 32'h13013019;
          16'h0b0f : blkif.rom_rdata <= 32'h23a02000;
          16'h0b10 : blkif.rom_rdata <= 32'h97500000;
          16'h0b11 : blkif.rom_rdata <= 32'h9380e03d;
          16'h0b12 : blkif.rom_rdata <= 32'h1301a00a;
          16'h0b13 : blkif.rom_rdata <= 32'h239d20fe;
          16'h0b14 : blkif.rom_rdata <= 32'h8391a0ff;
          16'h0b15 : blkif.rom_rdata <= 32'h930ea00a;
          16'h0b16 : blkif.rom_rdata <= 32'h130e3019;
          16'h0b17 : blkif.rom_rdata <= 32'h6384d101;
          16'h0b18 : blkif.rom_rdata <= 32'h6f20d030;
          16'h0b19 : blkif.rom_rdata <= 32'hb7000080;
          16'h0b1a : blkif.rom_rdata <= 32'h93804000;
          16'h0b1b : blkif.rom_rdata <= 32'h13014019;
          16'h0b1c : blkif.rom_rdata <= 32'h23a02000;
          16'h0b1d : blkif.rom_rdata <= 32'h97500000;
          16'h0b1e : blkif.rom_rdata <= 32'h9380a03a;
          16'h0b1f : blkif.rom_rdata <= 32'h37b1ffff;
          16'h0b20 : blkif.rom_rdata <= 32'h130101a0;
          16'h0b21 : blkif.rom_rdata <= 32'h239e20fe;
          16'h0b22 : blkif.rom_rdata <= 32'h8391c0ff;
          16'h0b23 : blkif.rom_rdata <= 32'hb7beffff;
          16'h0b24 : blkif.rom_rdata <= 32'h938e0ea0;
          16'h0b25 : blkif.rom_rdata <= 32'h130e4019;
          16'h0b26 : blkif.rom_rdata <= 32'h6384d101;
          16'h0b27 : blkif.rom_rdata <= 32'h6f20102d;
          16'h0b28 : blkif.rom_rdata <= 32'hb7000080;
          16'h0b29 : blkif.rom_rdata <= 32'h93804000;
          16'h0b2a : blkif.rom_rdata <= 32'h13016019;
          16'h0b2b : blkif.rom_rdata <= 32'h23a02000;
          16'h0b2c : blkif.rom_rdata <= 32'h97500000;
          16'h0b2d : blkif.rom_rdata <= 32'h9380e036;
          16'h0b2e : blkif.rom_rdata <= 32'h37a1ffff;
          16'h0b2f : blkif.rom_rdata <= 32'h1301a100;
          16'h0b30 : blkif.rom_rdata <= 32'h23902000;
          16'h0b31 : blkif.rom_rdata <= 32'h83910000;
          16'h0b32 : blkif.rom_rdata <= 32'hb7aeffff;
          16'h0b33 : blkif.rom_rdata <= 32'h938eae00;
          16'h0b34 : blkif.rom_rdata <= 32'h130e6019;
          16'h0b35 : blkif.rom_rdata <= 32'h6384d101;
          16'h0b36 : blkif.rom_rdata <= 32'h6f205029;
          16'h0b37 : blkif.rom_rdata <= 32'hb7000080;
          16'h0b38 : blkif.rom_rdata <= 32'h93804000;
          16'h0b39 : blkif.rom_rdata <= 32'h13017019;
          16'h0b3a : blkif.rom_rdata <= 32'h23a02000;
          16'h0b3b : blkif.rom_rdata <= 32'h97500000;
          16'h0b3c : blkif.rom_rdata <= 32'h93804033;
          16'h0b3d : blkif.rom_rdata <= 32'h37513412;
          16'h0b3e : blkif.rom_rdata <= 32'h13018167;
          16'h0b3f : blkif.rom_rdata <= 32'h138200fe;
          16'h0b40 : blkif.rom_rdata <= 32'h23102202;
          16'h0b41 : blkif.rom_rdata <= 32'h83910000;
          16'h0b42 : blkif.rom_rdata <= 32'hb75e0000;
          16'h0b43 : blkif.rom_rdata <= 32'h938e8e67;
          16'h0b44 : blkif.rom_rdata <= 32'h130e7019;
          16'h0b45 : blkif.rom_rdata <= 32'h6384d101;
          16'h0b46 : blkif.rom_rdata <= 32'h6f205025;
          16'h0b47 : blkif.rom_rdata <= 32'hb7000080;
          16'h0b48 : blkif.rom_rdata <= 32'h93804000;
          16'h0b49 : blkif.rom_rdata <= 32'h13018019;
          16'h0b4a : blkif.rom_rdata <= 32'h23a02000;
          16'h0b4b : blkif.rom_rdata <= 32'h97500000;
          16'h0b4c : blkif.rom_rdata <= 32'h9380402f;
          16'h0b4d : blkif.rom_rdata <= 32'h37310000;
          16'h0b4e : blkif.rom_rdata <= 32'h13018109;
          16'h0b4f : blkif.rom_rdata <= 32'h9380b0ff;
          16'h0b50 : blkif.rom_rdata <= 32'ha3932000;
          16'h0b51 : blkif.rom_rdata <= 32'h17520000;
          16'h0b52 : blkif.rom_rdata <= 32'h1302e22d;
          16'h0b53 : blkif.rom_rdata <= 32'h83110200;
          16'h0b54 : blkif.rom_rdata <= 32'hb73e0000;
          16'h0b55 : blkif.rom_rdata <= 32'h938e8e09;
          16'h0b56 : blkif.rom_rdata <= 32'h130e8019;
          16'h0b57 : blkif.rom_rdata <= 32'h6384d101;
          16'h0b58 : blkif.rom_rdata <= 32'h6f20d020;
          16'h0b59 : blkif.rom_rdata <= 32'h130e9019;
          16'h0b5a : blkif.rom_rdata <= 32'h13020000;
          16'h0b5b : blkif.rom_rdata <= 32'hb7d0ffff;
          16'h0b5c : blkif.rom_rdata <= 32'h9380d0cd;
          16'h0b5d : blkif.rom_rdata <= 32'h17510000;
          16'h0b5e : blkif.rom_rdata <= 32'h1301c129;
          16'h0b5f : blkif.rom_rdata <= 32'h23101100;
          16'h0b60 : blkif.rom_rdata <= 32'h83110100;
          16'h0b61 : blkif.rom_rdata <= 32'hb7deffff;
          16'h0b62 : blkif.rom_rdata <= 32'h938edecd;
          16'h0b63 : blkif.rom_rdata <= 32'h6384d101;
          16'h0b64 : blkif.rom_rdata <= 32'h6f20d01d;
          16'h0b65 : blkif.rom_rdata <= 32'h13021200;
          16'h0b66 : blkif.rom_rdata <= 32'h93022000;
          16'h0b67 : blkif.rom_rdata <= 32'he31852fc;
          16'h0b68 : blkif.rom_rdata <= 32'h130ee019;
          16'h0b69 : blkif.rom_rdata <= 32'h13020000;
          16'h0b6a : blkif.rom_rdata <= 32'hb7e0ffff;
          16'h0b6b : blkif.rom_rdata <= 32'h9380b0aa;
          16'h0b6c : blkif.rom_rdata <= 32'h13000000;
          16'h0b6d : blkif.rom_rdata <= 32'h13000000;
          16'h0b6e : blkif.rom_rdata <= 32'h17510000;
          16'h0b6f : blkif.rom_rdata <= 32'h13018125;
          16'h0b70 : blkif.rom_rdata <= 32'h23151100;
          16'h0b71 : blkif.rom_rdata <= 32'h8311a100;
          16'h0b72 : blkif.rom_rdata <= 32'hb7eeffff;
          16'h0b73 : blkif.rom_rdata <= 32'h938ebeaa;
          16'h0b74 : blkif.rom_rdata <= 32'h6384d101;
          16'h0b75 : blkif.rom_rdata <= 32'h6f209019;
          16'h0b76 : blkif.rom_rdata <= 32'h13021200;
          16'h0b77 : blkif.rom_rdata <= 32'h93022000;
          16'h0b78 : blkif.rom_rdata <= 32'he31452fc;
          16'h0b79 : blkif.rom_rdata <= 32'h130ef019;
          16'h0b7a : blkif.rom_rdata <= 32'h13020000;
          16'h0b7b : blkif.rom_rdata <= 32'h17510000;
          16'h0b7c : blkif.rom_rdata <= 32'h13014122;
          16'h0b7d : blkif.rom_rdata <= 32'hb7200000;
          16'h0b7e : blkif.rom_rdata <= 32'h93803023;
          16'h0b7f : blkif.rom_rdata <= 32'h23101100;
          16'h0b80 : blkif.rom_rdata <= 32'h83110100;
          16'h0b81 : blkif.rom_rdata <= 32'hb72e0000;
          16'h0b82 : blkif.rom_rdata <= 32'h938e3e23;
          16'h0b83 : blkif.rom_rdata <= 32'h6384d101;
          16'h0b84 : blkif.rom_rdata <= 32'h6f20d015;
          16'h0b85 : blkif.rom_rdata <= 32'h13021200;
          16'h0b86 : blkif.rom_rdata <= 32'h93022000;
          16'h0b87 : blkif.rom_rdata <= 32'he31852fc;
          16'h0b88 : blkif.rom_rdata <= 32'h130e301a;
          16'h0b89 : blkif.rom_rdata <= 32'h13020000;
          16'h0b8a : blkif.rom_rdata <= 32'h17510000;
          16'h0b8b : blkif.rom_rdata <= 32'h1301811e;
          16'h0b8c : blkif.rom_rdata <= 32'h13000000;
          16'h0b8d : blkif.rom_rdata <= 32'h93001001;
          16'h0b8e : blkif.rom_rdata <= 32'h13000000;
          16'h0b8f : blkif.rom_rdata <= 32'h23141100;
          16'h0b90 : blkif.rom_rdata <= 32'h83118100;
          16'h0b91 : blkif.rom_rdata <= 32'h930e1001;
          16'h0b92 : blkif.rom_rdata <= 32'h6384d101;
          16'h0b93 : blkif.rom_rdata <= 32'h6f201012;
          16'h0b94 : blkif.rom_rdata <= 32'h13021200;
          16'h0b95 : blkif.rom_rdata <= 32'h93022000;
          16'h0b96 : blkif.rom_rdata <= 32'he31852fc;
          16'h0b97 : blkif.rom_rdata <= 32'h130e401a;
          16'h0b98 : blkif.rom_rdata <= 32'h13020000;
          16'h0b99 : blkif.rom_rdata <= 32'h17510000;
          16'h0b9a : blkif.rom_rdata <= 32'h1301c11a;
          16'h0b9b : blkif.rom_rdata <= 32'h13000000;
          16'h0b9c : blkif.rom_rdata <= 32'h13000000;
          16'h0b9d : blkif.rom_rdata <= 32'hb7300000;
          16'h0b9e : blkif.rom_rdata <= 32'h93801000;
          16'h0b9f : blkif.rom_rdata <= 32'h23151100;
          16'h0ba0 : blkif.rom_rdata <= 32'h8311a100;
          16'h0ba1 : blkif.rom_rdata <= 32'hb73e0000;
          16'h0ba2 : blkif.rom_rdata <= 32'h938e1e00;
          16'h0ba3 : blkif.rom_rdata <= 32'h6384d101;
          16'h0ba4 : blkif.rom_rdata <= 32'h6f20d00d;
          16'h0ba5 : blkif.rom_rdata <= 32'h13021200;
          16'h0ba6 : blkif.rom_rdata <= 32'h93022000;
          16'h0ba7 : blkif.rom_rdata <= 32'he31452fc;
          16'h0ba8 : blkif.rom_rdata <= 32'h37c50000;
          16'h0ba9 : blkif.rom_rdata <= 32'h1305f5ee;
          16'h0baa : blkif.rom_rdata <= 32'h97550000;
          16'h0bab : blkif.rom_rdata <= 32'h93858516;
          16'h0bac : blkif.rom_rdata <= 32'h2393a500;
          16'h0bad : blkif.rom_rdata <= 32'hb7000080;
          16'h0bae : blkif.rom_rdata <= 32'h93804000;
          16'h0baf : blkif.rom_rdata <= 32'h1301501a;
          16'h0bb0 : blkif.rom_rdata <= 32'h23a02000;
          16'h0bb1 : blkif.rom_rdata <= 32'h93001000;
          16'h0bb2 : blkif.rom_rdata <= 32'h13010000;
          16'h0bb3 : blkif.rom_rdata <= 32'hb3912000;
          16'h0bb4 : blkif.rom_rdata <= 32'h930e1000;
          16'h0bb5 : blkif.rom_rdata <= 32'h130e501a;
          16'h0bb6 : blkif.rom_rdata <= 32'h6384d101;
          16'h0bb7 : blkif.rom_rdata <= 32'h6f201009;
          16'h0bb8 : blkif.rom_rdata <= 32'hb7000080;
          16'h0bb9 : blkif.rom_rdata <= 32'h93804000;
          16'h0bba : blkif.rom_rdata <= 32'h1301601a;
          16'h0bbb : blkif.rom_rdata <= 32'h23a02000;
          16'h0bbc : blkif.rom_rdata <= 32'h93001000;
          16'h0bbd : blkif.rom_rdata <= 32'h13011000;
          16'h0bbe : blkif.rom_rdata <= 32'hb3912000;
          16'h0bbf : blkif.rom_rdata <= 32'h930e2000;
          16'h0bc0 : blkif.rom_rdata <= 32'h130e601a;
          16'h0bc1 : blkif.rom_rdata <= 32'h6384d101;
          16'h0bc2 : blkif.rom_rdata <= 32'h6f205006;
          16'h0bc3 : blkif.rom_rdata <= 32'hb7000080;
          16'h0bc4 : blkif.rom_rdata <= 32'h93804000;
          16'h0bc5 : blkif.rom_rdata <= 32'h1301701a;
          16'h0bc6 : blkif.rom_rdata <= 32'h23a02000;
          16'h0bc7 : blkif.rom_rdata <= 32'h93001000;
          16'h0bc8 : blkif.rom_rdata <= 32'h13017000;
          16'h0bc9 : blkif.rom_rdata <= 32'hb3912000;
          16'h0bca : blkif.rom_rdata <= 32'h930e0008;
          16'h0bcb : blkif.rom_rdata <= 32'h130e701a;
          16'h0bcc : blkif.rom_rdata <= 32'h6384d101;
          16'h0bcd : blkif.rom_rdata <= 32'h6f209003;
          16'h0bce : blkif.rom_rdata <= 32'hb7000080;
          16'h0bcf : blkif.rom_rdata <= 32'h93804000;
          16'h0bd0 : blkif.rom_rdata <= 32'h1301a01a;
          16'h0bd1 : blkif.rom_rdata <= 32'h23a02000;
          16'h0bd2 : blkif.rom_rdata <= 32'h9300f0ff;
          16'h0bd3 : blkif.rom_rdata <= 32'h13010000;
          16'h0bd4 : blkif.rom_rdata <= 32'hb3912000;
          16'h0bd5 : blkif.rom_rdata <= 32'h930ef0ff;
          16'h0bd6 : blkif.rom_rdata <= 32'h130ea01a;
          16'h0bd7 : blkif.rom_rdata <= 32'h6384d101;
          16'h0bd8 : blkif.rom_rdata <= 32'h6f20d000;
          16'h0bd9 : blkif.rom_rdata <= 32'hb7000080;
          16'h0bda : blkif.rom_rdata <= 32'h93804000;
          16'h0bdb : blkif.rom_rdata <= 32'h1301e01a;
          16'h0bdc : blkif.rom_rdata <= 32'h23a02000;
          16'h0bdd : blkif.rom_rdata <= 32'h9300f0ff;
          16'h0bde : blkif.rom_rdata <= 32'h1301f001;
          16'h0bdf : blkif.rom_rdata <= 32'hb3912000;
          16'h0be0 : blkif.rom_rdata <= 32'hb70e0080;
          16'h0be1 : blkif.rom_rdata <= 32'h130ee01a;
          16'h0be2 : blkif.rom_rdata <= 32'h6384d101;
          16'h0be3 : blkif.rom_rdata <= 32'h6f20007e;
          16'h0be4 : blkif.rom_rdata <= 32'hb7000080;
          16'h0be5 : blkif.rom_rdata <= 32'h93804000;
          16'h0be6 : blkif.rom_rdata <= 32'h1301201b;
          16'h0be7 : blkif.rom_rdata <= 32'h23a02000;
          16'h0be8 : blkif.rom_rdata <= 32'hb7202121;
          16'h0be9 : blkif.rom_rdata <= 32'h93801012;
          16'h0bea : blkif.rom_rdata <= 32'h1301e000;
          16'h0beb : blkif.rom_rdata <= 32'hb3912000;
          16'h0bec : blkif.rom_rdata <= 32'hb74e4848;
          16'h0bed : blkif.rom_rdata <= 32'h130e201b;
          16'h0bee : blkif.rom_rdata <= 32'h6384d101;
          16'h0bef : blkif.rom_rdata <= 32'h6f20007b;
          16'h0bf0 : blkif.rom_rdata <= 32'hb7000080;
          16'h0bf1 : blkif.rom_rdata <= 32'h93804000;
          16'h0bf2 : blkif.rom_rdata <= 32'h1301301b;
          16'h0bf3 : blkif.rom_rdata <= 32'h23a02000;
          16'h0bf4 : blkif.rom_rdata <= 32'hb7202121;
          16'h0bf5 : blkif.rom_rdata <= 32'h93801012;
          16'h0bf6 : blkif.rom_rdata <= 32'h1301f001;
          16'h0bf7 : blkif.rom_rdata <= 32'hb3912000;
          16'h0bf8 : blkif.rom_rdata <= 32'hb70e0080;
          16'h0bf9 : blkif.rom_rdata <= 32'h130e301b;
          16'h0bfa : blkif.rom_rdata <= 32'h6384d101;
          16'h0bfb : blkif.rom_rdata <= 32'h6f200078;
          16'h0bfc : blkif.rom_rdata <= 32'hb7000080;
          16'h0bfd : blkif.rom_rdata <= 32'h93804000;
          16'h0bfe : blkif.rom_rdata <= 32'h1301401b;
          16'h0bff : blkif.rom_rdata <= 32'h23a02000;
          16'h0c00 : blkif.rom_rdata <= 32'hb7202121;
          16'h0c01 : blkif.rom_rdata <= 32'h93801012;
          16'h0c02 : blkif.rom_rdata <= 32'h130100fe;
          16'h0c03 : blkif.rom_rdata <= 32'hb3912000;
          16'h0c04 : blkif.rom_rdata <= 32'hb72e2121;
          16'h0c05 : blkif.rom_rdata <= 32'h938e1e12;
          16'h0c06 : blkif.rom_rdata <= 32'h130e401b;
          16'h0c07 : blkif.rom_rdata <= 32'h6384d101;
          16'h0c08 : blkif.rom_rdata <= 32'h6f20c074;
          16'h0c09 : blkif.rom_rdata <= 32'hb7000080;
          16'h0c0a : blkif.rom_rdata <= 32'h93804000;
          16'h0c0b : blkif.rom_rdata <= 32'h1301501b;
          16'h0c0c : blkif.rom_rdata <= 32'h23a02000;
          16'h0c0d : blkif.rom_rdata <= 32'hb7202121;
          16'h0c0e : blkif.rom_rdata <= 32'h93801012;
          16'h0c0f : blkif.rom_rdata <= 32'h130110fe;
          16'h0c10 : blkif.rom_rdata <= 32'hb3912000;
          16'h0c11 : blkif.rom_rdata <= 32'hb74e4242;
          16'h0c12 : blkif.rom_rdata <= 32'h938e2e24;
          16'h0c13 : blkif.rom_rdata <= 32'h130e501b;
          16'h0c14 : blkif.rom_rdata <= 32'h6384d101;
          16'h0c15 : blkif.rom_rdata <= 32'h6f208071;
          16'h0c16 : blkif.rom_rdata <= 32'hb7000080;
          16'h0c17 : blkif.rom_rdata <= 32'h93804000;
          16'h0c18 : blkif.rom_rdata <= 32'h1301601b;
          16'h0c19 : blkif.rom_rdata <= 32'h23a02000;
          16'h0c1a : blkif.rom_rdata <= 32'hb7202121;
          16'h0c1b : blkif.rom_rdata <= 32'h93801012;
          16'h0c1c : blkif.rom_rdata <= 32'h130170fe;
          16'h0c1d : blkif.rom_rdata <= 32'hb3912000;
          16'h0c1e : blkif.rom_rdata <= 32'hb79e9090;
          16'h0c1f : blkif.rom_rdata <= 32'h938e0e08;
          16'h0c20 : blkif.rom_rdata <= 32'h130e601b;
          16'h0c21 : blkif.rom_rdata <= 32'h6384d101;
          16'h0c22 : blkif.rom_rdata <= 32'h6f20406e;
          16'h0c23 : blkif.rom_rdata <= 32'hb7000080;
          16'h0c24 : blkif.rom_rdata <= 32'h93804000;
          16'h0c25 : blkif.rom_rdata <= 32'h1301701b;
          16'h0c26 : blkif.rom_rdata <= 32'h23a02000;
          16'h0c27 : blkif.rom_rdata <= 32'hb7202121;
          16'h0c28 : blkif.rom_rdata <= 32'h93801012;
          16'h0c29 : blkif.rom_rdata <= 32'h1301e0fe;
          16'h0c2a : blkif.rom_rdata <= 32'hb3912000;
          16'h0c2b : blkif.rom_rdata <= 32'hb74e4848;
          16'h0c2c : blkif.rom_rdata <= 32'h130e701b;
          16'h0c2d : blkif.rom_rdata <= 32'h6384d101;
          16'h0c2e : blkif.rom_rdata <= 32'h6f20406b;
          16'h0c2f : blkif.rom_rdata <= 32'hb7000080;
          16'h0c30 : blkif.rom_rdata <= 32'h93804000;
          16'h0c31 : blkif.rom_rdata <= 32'h1301801b;
          16'h0c32 : blkif.rom_rdata <= 32'h23a02000;
          16'h0c33 : blkif.rom_rdata <= 32'hb7202121;
          16'h0c34 : blkif.rom_rdata <= 32'h93800012;
          16'h0c35 : blkif.rom_rdata <= 32'h1301f0ff;
          16'h0c36 : blkif.rom_rdata <= 32'hb3912000;
          16'h0c37 : blkif.rom_rdata <= 32'h930e0000;
          16'h0c38 : blkif.rom_rdata <= 32'h130e801b;
          16'h0c39 : blkif.rom_rdata <= 32'h6384d101;
          16'h0c3a : blkif.rom_rdata <= 32'h6f204068;
          16'h0c3b : blkif.rom_rdata <= 32'hb7000080;
          16'h0c3c : blkif.rom_rdata <= 32'h93804000;
          16'h0c3d : blkif.rom_rdata <= 32'h1301901b;
          16'h0c3e : blkif.rom_rdata <= 32'h23a02000;
          16'h0c3f : blkif.rom_rdata <= 32'h93001000;
          16'h0c40 : blkif.rom_rdata <= 32'h13017000;
          16'h0c41 : blkif.rom_rdata <= 32'hb3902000;
          16'h0c42 : blkif.rom_rdata <= 32'h930e0008;
          16'h0c43 : blkif.rom_rdata <= 32'h130e901b;
          16'h0c44 : blkif.rom_rdata <= 32'h6384d001;
          16'h0c45 : blkif.rom_rdata <= 32'h6f208065;
          16'h0c46 : blkif.rom_rdata <= 32'hb7000080;
          16'h0c47 : blkif.rom_rdata <= 32'h93804000;
          16'h0c48 : blkif.rom_rdata <= 32'h1301a01b;
          16'h0c49 : blkif.rom_rdata <= 32'h23a02000;
          16'h0c4a : blkif.rom_rdata <= 32'h93001000;
          16'h0c4b : blkif.rom_rdata <= 32'h1301e000;
          16'h0c4c : blkif.rom_rdata <= 32'h33912000;
          16'h0c4d : blkif.rom_rdata <= 32'hb74e0000;
          16'h0c4e : blkif.rom_rdata <= 32'h130ea01b;
          16'h0c4f : blkif.rom_rdata <= 32'h6304d101;
          16'h0c50 : blkif.rom_rdata <= 32'h6f20c062;
          16'h0c51 : blkif.rom_rdata <= 32'hb7000080;
          16'h0c52 : blkif.rom_rdata <= 32'h93804000;
          16'h0c53 : blkif.rom_rdata <= 32'h1301b01b;
          16'h0c54 : blkif.rom_rdata <= 32'h23a02000;
          16'h0c55 : blkif.rom_rdata <= 32'h93003000;
          16'h0c56 : blkif.rom_rdata <= 32'hb3901000;
          16'h0c57 : blkif.rom_rdata <= 32'h930e8001;
          16'h0c58 : blkif.rom_rdata <= 32'h130eb01b;
          16'h0c59 : blkif.rom_rdata <= 32'h6384d001;
          16'h0c5a : blkif.rom_rdata <= 32'h6f204060;
          16'h0c5b : blkif.rom_rdata <= 32'hb7000080;
          16'h0c5c : blkif.rom_rdata <= 32'h93804000;
          16'h0c5d : blkif.rom_rdata <= 32'h1301c01b;
          16'h0c5e : blkif.rom_rdata <= 32'h23a02000;
          16'h0c5f : blkif.rom_rdata <= 32'h13020000;
          16'h0c60 : blkif.rom_rdata <= 32'h93001000;
          16'h0c61 : blkif.rom_rdata <= 32'h13017000;
          16'h0c62 : blkif.rom_rdata <= 32'hb3912000;
          16'h0c63 : blkif.rom_rdata <= 32'h13830100;
          16'h0c64 : blkif.rom_rdata <= 32'h13021200;
          16'h0c65 : blkif.rom_rdata <= 32'h93022000;
          16'h0c66 : blkif.rom_rdata <= 32'he31452fe;
          16'h0c67 : blkif.rom_rdata <= 32'h930e0008;
          16'h0c68 : blkif.rom_rdata <= 32'h130ec01b;
          16'h0c69 : blkif.rom_rdata <= 32'h6304d301;
          16'h0c6a : blkif.rom_rdata <= 32'h6f20405c;
          16'h0c6b : blkif.rom_rdata <= 32'hb7000080;
          16'h0c6c : blkif.rom_rdata <= 32'h93804000;
          16'h0c6d : blkif.rom_rdata <= 32'h1301d01b;
          16'h0c6e : blkif.rom_rdata <= 32'h23a02000;
          16'h0c6f : blkif.rom_rdata <= 32'h13020000;
          16'h0c70 : blkif.rom_rdata <= 32'h93001000;
          16'h0c71 : blkif.rom_rdata <= 32'h1301e000;
          16'h0c72 : blkif.rom_rdata <= 32'hb3912000;
          16'h0c73 : blkif.rom_rdata <= 32'h13000000;
          16'h0c74 : blkif.rom_rdata <= 32'h13830100;
          16'h0c75 : blkif.rom_rdata <= 32'h13021200;
          16'h0c76 : blkif.rom_rdata <= 32'h93022000;
          16'h0c77 : blkif.rom_rdata <= 32'he31252fe;
          16'h0c78 : blkif.rom_rdata <= 32'hb74e0000;
          16'h0c79 : blkif.rom_rdata <= 32'h130ed01b;
          16'h0c7a : blkif.rom_rdata <= 32'h6304d301;
          16'h0c7b : blkif.rom_rdata <= 32'h6f200058;
          16'h0c7c : blkif.rom_rdata <= 32'hb7000080;
          16'h0c7d : blkif.rom_rdata <= 32'h93804000;
          16'h0c7e : blkif.rom_rdata <= 32'h1301e01b;
          16'h0c7f : blkif.rom_rdata <= 32'h23a02000;
          16'h0c80 : blkif.rom_rdata <= 32'h13020000;
          16'h0c81 : blkif.rom_rdata <= 32'h93001000;
          16'h0c82 : blkif.rom_rdata <= 32'h1301f001;
          16'h0c83 : blkif.rom_rdata <= 32'hb3912000;
          16'h0c84 : blkif.rom_rdata <= 32'h13000000;
          16'h0c85 : blkif.rom_rdata <= 32'h13000000;
          16'h0c86 : blkif.rom_rdata <= 32'h13830100;
          16'h0c87 : blkif.rom_rdata <= 32'h13021200;
          16'h0c88 : blkif.rom_rdata <= 32'h93022000;
          16'h0c89 : blkif.rom_rdata <= 32'he31052fe;
          16'h0c8a : blkif.rom_rdata <= 32'hb70e0080;
          16'h0c8b : blkif.rom_rdata <= 32'h130ee01b;
          16'h0c8c : blkif.rom_rdata <= 32'h6304d301;
          16'h0c8d : blkif.rom_rdata <= 32'h6f208053;
          16'h0c8e : blkif.rom_rdata <= 32'hb7000080;
          16'h0c8f : blkif.rom_rdata <= 32'h93804000;
          16'h0c90 : blkif.rom_rdata <= 32'h1301f01b;
          16'h0c91 : blkif.rom_rdata <= 32'h23a02000;
          16'h0c92 : blkif.rom_rdata <= 32'h13020000;
          16'h0c93 : blkif.rom_rdata <= 32'h93001000;
          16'h0c94 : blkif.rom_rdata <= 32'h13017000;
          16'h0c95 : blkif.rom_rdata <= 32'hb3912000;
          16'h0c96 : blkif.rom_rdata <= 32'h13021200;
          16'h0c97 : blkif.rom_rdata <= 32'h93022000;
          16'h0c98 : blkif.rom_rdata <= 32'he31652fe;
          16'h0c99 : blkif.rom_rdata <= 32'h930e0008;
          16'h0c9a : blkif.rom_rdata <= 32'h130ef01b;
          16'h0c9b : blkif.rom_rdata <= 32'h6384d101;
          16'h0c9c : blkif.rom_rdata <= 32'h6f20c04f;
          16'h0c9d : blkif.rom_rdata <= 32'hb7000080;
          16'h0c9e : blkif.rom_rdata <= 32'h93804000;
          16'h0c9f : blkif.rom_rdata <= 32'h1301401c;
          16'h0ca0 : blkif.rom_rdata <= 32'h23a02000;
          16'h0ca1 : blkif.rom_rdata <= 32'h13020000;
          16'h0ca2 : blkif.rom_rdata <= 32'h93001000;
          16'h0ca3 : blkif.rom_rdata <= 32'h13000000;
          16'h0ca4 : blkif.rom_rdata <= 32'h13000000;
          16'h0ca5 : blkif.rom_rdata <= 32'h1301f001;
          16'h0ca6 : blkif.rom_rdata <= 32'hb3912000;
          16'h0ca7 : blkif.rom_rdata <= 32'h13021200;
          16'h0ca8 : blkif.rom_rdata <= 32'h93022000;
          16'h0ca9 : blkif.rom_rdata <= 32'he31252fe;
          16'h0caa : blkif.rom_rdata <= 32'hb70e0080;
          16'h0cab : blkif.rom_rdata <= 32'h130e401c;
          16'h0cac : blkif.rom_rdata <= 32'h6384d101;
          16'h0cad : blkif.rom_rdata <= 32'h6f20804b;
          16'h0cae : blkif.rom_rdata <= 32'hb7000080;
          16'h0caf : blkif.rom_rdata <= 32'h93804000;
          16'h0cb0 : blkif.rom_rdata <= 32'h1301501c;
          16'h0cb1 : blkif.rom_rdata <= 32'h23a02000;
          16'h0cb2 : blkif.rom_rdata <= 32'h13020000;
          16'h0cb3 : blkif.rom_rdata <= 32'h13017000;
          16'h0cb4 : blkif.rom_rdata <= 32'h93001000;
          16'h0cb5 : blkif.rom_rdata <= 32'hb3912000;
          16'h0cb6 : blkif.rom_rdata <= 32'h13021200;
          16'h0cb7 : blkif.rom_rdata <= 32'h93022000;
          16'h0cb8 : blkif.rom_rdata <= 32'he31652fe;
          16'h0cb9 : blkif.rom_rdata <= 32'h930e0008;
          16'h0cba : blkif.rom_rdata <= 32'h130e501c;
          16'h0cbb : blkif.rom_rdata <= 32'h6384d101;
          16'h0cbc : blkif.rom_rdata <= 32'h6f20c047;
          16'h0cbd : blkif.rom_rdata <= 32'hb7000080;
          16'h0cbe : blkif.rom_rdata <= 32'h93804000;
          16'h0cbf : blkif.rom_rdata <= 32'h1301a01c;
          16'h0cc0 : blkif.rom_rdata <= 32'h23a02000;
          16'h0cc1 : blkif.rom_rdata <= 32'h13020000;
          16'h0cc2 : blkif.rom_rdata <= 32'h1301f001;
          16'h0cc3 : blkif.rom_rdata <= 32'h13000000;
          16'h0cc4 : blkif.rom_rdata <= 32'h13000000;
          16'h0cc5 : blkif.rom_rdata <= 32'h93001000;
          16'h0cc6 : blkif.rom_rdata <= 32'hb3912000;
          16'h0cc7 : blkif.rom_rdata <= 32'h13021200;
          16'h0cc8 : blkif.rom_rdata <= 32'h93022000;
          16'h0cc9 : blkif.rom_rdata <= 32'he31252fe;
          16'h0cca : blkif.rom_rdata <= 32'hb70e0080;
          16'h0ccb : blkif.rom_rdata <= 32'h130ea01c;
          16'h0ccc : blkif.rom_rdata <= 32'h6384d101;
          16'h0ccd : blkif.rom_rdata <= 32'h6f208043;
          16'h0cce : blkif.rom_rdata <= 32'hb7000080;
          16'h0ccf : blkif.rom_rdata <= 32'h93804000;
          16'h0cd0 : blkif.rom_rdata <= 32'h1301b01c;
          16'h0cd1 : blkif.rom_rdata <= 32'h23a02000;
          16'h0cd2 : blkif.rom_rdata <= 32'h9300f000;
          16'h0cd3 : blkif.rom_rdata <= 32'h33111000;
          16'h0cd4 : blkif.rom_rdata <= 32'h930e0000;
          16'h0cd5 : blkif.rom_rdata <= 32'h130eb01c;
          16'h0cd6 : blkif.rom_rdata <= 32'h6304d101;
          16'h0cd7 : blkif.rom_rdata <= 32'h6f200041;
          16'h0cd8 : blkif.rom_rdata <= 32'hb7000080;
          16'h0cd9 : blkif.rom_rdata <= 32'h93804000;
          16'h0cda : blkif.rom_rdata <= 32'h1301c01c;
          16'h0cdb : blkif.rom_rdata <= 32'h23a02000;
          16'h0cdc : blkif.rom_rdata <= 32'h93000002;
          16'h0cdd : blkif.rom_rdata <= 32'h33910000;
          16'h0cde : blkif.rom_rdata <= 32'h930e0002;
          16'h0cdf : blkif.rom_rdata <= 32'h130ec01c;
          16'h0ce0 : blkif.rom_rdata <= 32'h6304d101;
          16'h0ce1 : blkif.rom_rdata <= 32'h6f20803e;
          16'h0ce2 : blkif.rom_rdata <= 32'hb7000080;
          16'h0ce3 : blkif.rom_rdata <= 32'h93804000;
          16'h0ce4 : blkif.rom_rdata <= 32'h1301d01c;
          16'h0ce5 : blkif.rom_rdata <= 32'h23a02000;
          16'h0ce6 : blkif.rom_rdata <= 32'hb3100000;
          16'h0ce7 : blkif.rom_rdata <= 32'h930e0000;
          16'h0ce8 : blkif.rom_rdata <= 32'h130ed01c;
          16'h0ce9 : blkif.rom_rdata <= 32'h6384d001;
          16'h0cea : blkif.rom_rdata <= 32'h6f20403c;
          16'h0ceb : blkif.rom_rdata <= 32'hb7000080;
          16'h0cec : blkif.rom_rdata <= 32'h93804000;
          16'h0ced : blkif.rom_rdata <= 32'h1301e01c;
          16'h0cee : blkif.rom_rdata <= 32'h23a02000;
          16'h0cef : blkif.rom_rdata <= 32'h93000040;
          16'h0cf0 : blkif.rom_rdata <= 32'h37110000;
          16'h0cf1 : blkif.rom_rdata <= 32'h13010180;
          16'h0cf2 : blkif.rom_rdata <= 32'h33902000;
          16'h0cf3 : blkif.rom_rdata <= 32'h930e0000;
          16'h0cf4 : blkif.rom_rdata <= 32'h130ee01c;
          16'h0cf5 : blkif.rom_rdata <= 32'h6304d001;
          16'h0cf6 : blkif.rom_rdata <= 32'h6f204039;
          16'h0cf7 : blkif.rom_rdata <= 32'hb7000080;
          16'h0cf8 : blkif.rom_rdata <= 32'h93804000;
          16'h0cf9 : blkif.rom_rdata <= 32'h1301f01c;
          16'h0cfa : blkif.rom_rdata <= 32'h23a02000;
          16'h0cfb : blkif.rom_rdata <= 32'h93001000;
          16'h0cfc : blkif.rom_rdata <= 32'h93910000;
          16'h0cfd : blkif.rom_rdata <= 32'h930e1000;
          16'h0cfe : blkif.rom_rdata <= 32'h130ef01c;
          16'h0cff : blkif.rom_rdata <= 32'h6384d101;
          16'h0d00 : blkif.rom_rdata <= 32'h6f20c036;
          16'h0d01 : blkif.rom_rdata <= 32'hb7000080;
          16'h0d02 : blkif.rom_rdata <= 32'h93804000;
          16'h0d03 : blkif.rom_rdata <= 32'h1301001d;
          16'h0d04 : blkif.rom_rdata <= 32'h23a02000;
          16'h0d05 : blkif.rom_rdata <= 32'h93001000;
          16'h0d06 : blkif.rom_rdata <= 32'h93911000;
          16'h0d07 : blkif.rom_rdata <= 32'h930e2000;
          16'h0d08 : blkif.rom_rdata <= 32'h130e001d;
          16'h0d09 : blkif.rom_rdata <= 32'h6384d101;
          16'h0d0a : blkif.rom_rdata <= 32'h6f204034;
          16'h0d0b : blkif.rom_rdata <= 32'hb7000080;
          16'h0d0c : blkif.rom_rdata <= 32'h93804000;
          16'h0d0d : blkif.rom_rdata <= 32'h1301301d;
          16'h0d0e : blkif.rom_rdata <= 32'h23a02000;
          16'h0d0f : blkif.rom_rdata <= 32'h93001000;
          16'h0d10 : blkif.rom_rdata <= 32'h9391f001;
          16'h0d11 : blkif.rom_rdata <= 32'hb70e0080;
          16'h0d12 : blkif.rom_rdata <= 32'h130e301d;
          16'h0d13 : blkif.rom_rdata <= 32'h6384d101;
          16'h0d14 : blkif.rom_rdata <= 32'h6f20c031;
          16'h0d15 : blkif.rom_rdata <= 32'hb7000080;
          16'h0d16 : blkif.rom_rdata <= 32'h93804000;
          16'h0d17 : blkif.rom_rdata <= 32'h1301401d;
          16'h0d18 : blkif.rom_rdata <= 32'h23a02000;
          16'h0d19 : blkif.rom_rdata <= 32'h9300f0ff;
          16'h0d1a : blkif.rom_rdata <= 32'h93910000;
          16'h0d1b : blkif.rom_rdata <= 32'h930ef0ff;
          16'h0d1c : blkif.rom_rdata <= 32'h130e401d;
          16'h0d1d : blkif.rom_rdata <= 32'h6384d101;
          16'h0d1e : blkif.rom_rdata <= 32'h6f20402f;
          16'h0d1f : blkif.rom_rdata <= 32'hb7000080;
          16'h0d20 : blkif.rom_rdata <= 32'h93804000;
          16'h0d21 : blkif.rom_rdata <= 32'h1301801d;
          16'h0d22 : blkif.rom_rdata <= 32'h23a02000;
          16'h0d23 : blkif.rom_rdata <= 32'h9300f0ff;
          16'h0d24 : blkif.rom_rdata <= 32'h9391f001;
          16'h0d25 : blkif.rom_rdata <= 32'hb70e0080;
          16'h0d26 : blkif.rom_rdata <= 32'h130e801d;
          16'h0d27 : blkif.rom_rdata <= 32'h6384d101;
          16'h0d28 : blkif.rom_rdata <= 32'h6f20c02c;
          16'h0d29 : blkif.rom_rdata <= 32'hb7000080;
          16'h0d2a : blkif.rom_rdata <= 32'h93804000;
          16'h0d2b : blkif.rom_rdata <= 32'h1301901d;
          16'h0d2c : blkif.rom_rdata <= 32'h23a02000;
          16'h0d2d : blkif.rom_rdata <= 32'hb7202121;
          16'h0d2e : blkif.rom_rdata <= 32'h93801012;
          16'h0d2f : blkif.rom_rdata <= 32'h93910000;
          16'h0d30 : blkif.rom_rdata <= 32'hb72e2121;
          16'h0d31 : blkif.rom_rdata <= 32'h938e1e12;
          16'h0d32 : blkif.rom_rdata <= 32'h130e901d;
          16'h0d33 : blkif.rom_rdata <= 32'h6384d101;
          16'h0d34 : blkif.rom_rdata <= 32'h6f20c029;
          16'h0d35 : blkif.rom_rdata <= 32'hb7000080;
          16'h0d36 : blkif.rom_rdata <= 32'h93804000;
          16'h0d37 : blkif.rom_rdata <= 32'h1301c01d;
          16'h0d38 : blkif.rom_rdata <= 32'h23a02000;
          16'h0d39 : blkif.rom_rdata <= 32'hb7202121;
          16'h0d3a : blkif.rom_rdata <= 32'h93801012;
          16'h0d3b : blkif.rom_rdata <= 32'h9391e000;
          16'h0d3c : blkif.rom_rdata <= 32'hb74e4848;
          16'h0d3d : blkif.rom_rdata <= 32'h130ec01d;
          16'h0d3e : blkif.rom_rdata <= 32'h6384d101;
          16'h0d3f : blkif.rom_rdata <= 32'h6f200027;
          16'h0d40 : blkif.rom_rdata <= 32'hb7000080;
          16'h0d41 : blkif.rom_rdata <= 32'h93804000;
          16'h0d42 : blkif.rom_rdata <= 32'h1301d01d;
          16'h0d43 : blkif.rom_rdata <= 32'h23a02000;
          16'h0d44 : blkif.rom_rdata <= 32'hb7202121;
          16'h0d45 : blkif.rom_rdata <= 32'h93801012;
          16'h0d46 : blkif.rom_rdata <= 32'h9391f001;
          16'h0d47 : blkif.rom_rdata <= 32'hb70e0080;
          16'h0d48 : blkif.rom_rdata <= 32'h130ed01d;
          16'h0d49 : blkif.rom_rdata <= 32'h6384d101;
          16'h0d4a : blkif.rom_rdata <= 32'h6f204024;
          16'h0d4b : blkif.rom_rdata <= 32'hb7000080;
          16'h0d4c : blkif.rom_rdata <= 32'h93804000;
          16'h0d4d : blkif.rom_rdata <= 32'h1301e01d;
          16'h0d4e : blkif.rom_rdata <= 32'h23a02000;
          16'h0d4f : blkif.rom_rdata <= 32'h93001000;
          16'h0d50 : blkif.rom_rdata <= 32'h93907000;
          16'h0d51 : blkif.rom_rdata <= 32'h930e0008;
          16'h0d52 : blkif.rom_rdata <= 32'h130ee01d;
          16'h0d53 : blkif.rom_rdata <= 32'h6384d001;
          16'h0d54 : blkif.rom_rdata <= 32'h6f20c021;
          16'h0d55 : blkif.rom_rdata <= 32'hb7000080;
          16'h0d56 : blkif.rom_rdata <= 32'h93804000;
          16'h0d57 : blkif.rom_rdata <= 32'h1301101e;
          16'h0d58 : blkif.rom_rdata <= 32'h23a02000;
          16'h0d59 : blkif.rom_rdata <= 32'h13020000;
          16'h0d5a : blkif.rom_rdata <= 32'h93001000;
          16'h0d5b : blkif.rom_rdata <= 32'h9391f001;
          16'h0d5c : blkif.rom_rdata <= 32'h13000000;
          16'h0d5d : blkif.rom_rdata <= 32'h13000000;
          16'h0d5e : blkif.rom_rdata <= 32'h13830100;
          16'h0d5f : blkif.rom_rdata <= 32'h13021200;
          16'h0d60 : blkif.rom_rdata <= 32'h93022000;
          16'h0d61 : blkif.rom_rdata <= 32'he31252fe;
          16'h0d62 : blkif.rom_rdata <= 32'hb70e0080;
          16'h0d63 : blkif.rom_rdata <= 32'h130e101e;
          16'h0d64 : blkif.rom_rdata <= 32'h6304d301;
          16'h0d65 : blkif.rom_rdata <= 32'h6f20801d;
          16'h0d66 : blkif.rom_rdata <= 32'hb7000080;
          16'h0d67 : blkif.rom_rdata <= 32'h93804000;
          16'h0d68 : blkif.rom_rdata <= 32'h1301201e;
          16'h0d69 : blkif.rom_rdata <= 32'h23a02000;
          16'h0d6a : blkif.rom_rdata <= 32'h13020000;
          16'h0d6b : blkif.rom_rdata <= 32'h93001000;
          16'h0d6c : blkif.rom_rdata <= 32'h93917000;
          16'h0d6d : blkif.rom_rdata <= 32'h13021200;
          16'h0d6e : blkif.rom_rdata <= 32'h93022000;
          16'h0d6f : blkif.rom_rdata <= 32'he31852fe;
          16'h0d70 : blkif.rom_rdata <= 32'h930e0008;
          16'h0d71 : blkif.rom_rdata <= 32'h130e201e;
          16'h0d72 : blkif.rom_rdata <= 32'h6384d101;
          16'h0d73 : blkif.rom_rdata <= 32'h6f20001a;
          16'h0d74 : blkif.rom_rdata <= 32'hb7000080;
          16'h0d75 : blkif.rom_rdata <= 32'h93804000;
          16'h0d76 : blkif.rom_rdata <= 32'h1301301e;
          16'h0d77 : blkif.rom_rdata <= 32'h23a02000;
          16'h0d78 : blkif.rom_rdata <= 32'h13020000;
          16'h0d79 : blkif.rom_rdata <= 32'h93001000;
          16'h0d7a : blkif.rom_rdata <= 32'h13000000;
          16'h0d7b : blkif.rom_rdata <= 32'h9391e000;
          16'h0d7c : blkif.rom_rdata <= 32'h13021200;
          16'h0d7d : blkif.rom_rdata <= 32'h93022000;
          16'h0d7e : blkif.rom_rdata <= 32'he31652fe;
          16'h0d7f : blkif.rom_rdata <= 32'hb74e0000;
          16'h0d80 : blkif.rom_rdata <= 32'h130e301e;
          16'h0d81 : blkif.rom_rdata <= 32'h6384d101;
          16'h0d82 : blkif.rom_rdata <= 32'h6f204016;
          16'h0d83 : blkif.rom_rdata <= 32'hb7000080;
          16'h0d84 : blkif.rom_rdata <= 32'h93804000;
          16'h0d85 : blkif.rom_rdata <= 32'h1301501e;
          16'h0d86 : blkif.rom_rdata <= 32'h23a02000;
          16'h0d87 : blkif.rom_rdata <= 32'h9310f001;
          16'h0d88 : blkif.rom_rdata <= 32'h930e0000;
          16'h0d89 : blkif.rom_rdata <= 32'h130e501e;
          16'h0d8a : blkif.rom_rdata <= 32'h6384d001;
          16'h0d8b : blkif.rom_rdata <= 32'h6f200014;
          16'h0d8c : blkif.rom_rdata <= 32'hb7000080;
          16'h0d8d : blkif.rom_rdata <= 32'h93804000;
          16'h0d8e : blkif.rom_rdata <= 32'h1301601e;
          16'h0d8f : blkif.rom_rdata <= 32'h23a02000;
          16'h0d90 : blkif.rom_rdata <= 32'h93001002;
          16'h0d91 : blkif.rom_rdata <= 32'h13904001;
          16'h0d92 : blkif.rom_rdata <= 32'h930e0000;
          16'h0d93 : blkif.rom_rdata <= 32'h130e601e;
          16'h0d94 : blkif.rom_rdata <= 32'h6304d001;
          16'h0d95 : blkif.rom_rdata <= 32'h6f208011;
          16'h0d96 : blkif.rom_rdata <= 32'hb7000080;
          16'h0d97 : blkif.rom_rdata <= 32'h93804000;
          16'h0d98 : blkif.rom_rdata <= 32'h1301701e;
          16'h0d99 : blkif.rom_rdata <= 32'h23a02000;
          16'h0d9a : blkif.rom_rdata <= 32'h93000000;
          16'h0d9b : blkif.rom_rdata <= 32'h13010000;
          16'h0d9c : blkif.rom_rdata <= 32'hb3a12000;
          16'h0d9d : blkif.rom_rdata <= 32'h930e0000;
          16'h0d9e : blkif.rom_rdata <= 32'h130e701e;
          16'h0d9f : blkif.rom_rdata <= 32'h6384d101;
          16'h0da0 : blkif.rom_rdata <= 32'h6f20c00e;
          16'h0da1 : blkif.rom_rdata <= 32'hb7000080;
          16'h0da2 : blkif.rom_rdata <= 32'h93804000;
          16'h0da3 : blkif.rom_rdata <= 32'h1301d01e;
          16'h0da4 : blkif.rom_rdata <= 32'h23a02000;
          16'h0da5 : blkif.rom_rdata <= 32'hb7000080;
          16'h0da6 : blkif.rom_rdata <= 32'h3781ffff;
          16'h0da7 : blkif.rom_rdata <= 32'hb3a12000;
          16'h0da8 : blkif.rom_rdata <= 32'h930e1000;
          16'h0da9 : blkif.rom_rdata <= 32'h130ed01e;
          16'h0daa : blkif.rom_rdata <= 32'h6384d101;
          16'h0dab : blkif.rom_rdata <= 32'h6f20000c;
          16'h0dac : blkif.rom_rdata <= 32'hb7000080;
          16'h0dad : blkif.rom_rdata <= 32'h93804000;
          16'h0dae : blkif.rom_rdata <= 32'h1301301f;
          16'h0daf : blkif.rom_rdata <= 32'h23a02000;
          16'h0db0 : blkif.rom_rdata <= 32'h93000000;
          16'h0db1 : blkif.rom_rdata <= 32'h1301f0ff;
          16'h0db2 : blkif.rom_rdata <= 32'hb3a12000;
          16'h0db3 : blkif.rom_rdata <= 32'h930e0000;
          16'h0db4 : blkif.rom_rdata <= 32'h130e301f;
          16'h0db5 : blkif.rom_rdata <= 32'h6384d101;
          16'h0db6 : blkif.rom_rdata <= 32'h6f204009;
          16'h0db7 : blkif.rom_rdata <= 32'hb7000080;
          16'h0db8 : blkif.rom_rdata <= 32'h93804000;
          16'h0db9 : blkif.rom_rdata <= 32'h1301501f;
          16'h0dba : blkif.rom_rdata <= 32'h23a02000;
          16'h0dbb : blkif.rom_rdata <= 32'h9300f0ff;
          16'h0dbc : blkif.rom_rdata <= 32'h1301f0ff;
          16'h0dbd : blkif.rom_rdata <= 32'hb3a12000;
          16'h0dbe : blkif.rom_rdata <= 32'h930e0000;
          16'h0dbf : blkif.rom_rdata <= 32'h130e501f;
          16'h0dc0 : blkif.rom_rdata <= 32'h6384d101;
          16'h0dc1 : blkif.rom_rdata <= 32'h6f208006;
          16'h0dc2 : blkif.rom_rdata <= 32'hb7000080;
          16'h0dc3 : blkif.rom_rdata <= 32'h93804000;
          16'h0dc4 : blkif.rom_rdata <= 32'h1301601f;
          16'h0dc5 : blkif.rom_rdata <= 32'h23a02000;
          16'h0dc6 : blkif.rom_rdata <= 32'h9300e000;
          16'h0dc7 : blkif.rom_rdata <= 32'h1301d000;
          16'h0dc8 : blkif.rom_rdata <= 32'hb3a02000;
          16'h0dc9 : blkif.rom_rdata <= 32'h930e0000;
          16'h0dca : blkif.rom_rdata <= 32'h130e601f;
          16'h0dcb : blkif.rom_rdata <= 32'h6384d001;
          16'h0dcc : blkif.rom_rdata <= 32'h6f20c003;
          16'h0dcd : blkif.rom_rdata <= 32'hb7000080;
          16'h0dce : blkif.rom_rdata <= 32'h93804000;
          16'h0dcf : blkif.rom_rdata <= 32'h1301701f;
          16'h0dd0 : blkif.rom_rdata <= 32'h23a02000;
          16'h0dd1 : blkif.rom_rdata <= 32'h9300b000;
          16'h0dd2 : blkif.rom_rdata <= 32'h1301d000;
          16'h0dd3 : blkif.rom_rdata <= 32'h33a12000;
          16'h0dd4 : blkif.rom_rdata <= 32'h930e1000;
          16'h0dd5 : blkif.rom_rdata <= 32'h130e701f;
          16'h0dd6 : blkif.rom_rdata <= 32'h6304d101;
          16'h0dd7 : blkif.rom_rdata <= 32'h6f200001;
          16'h0dd8 : blkif.rom_rdata <= 32'hb7000080;
          16'h0dd9 : blkif.rom_rdata <= 32'h93804000;
          16'h0dda : blkif.rom_rdata <= 32'h1301801f;
          16'h0ddb : blkif.rom_rdata <= 32'h23a02000;
          16'h0ddc : blkif.rom_rdata <= 32'h9300d000;
          16'h0ddd : blkif.rom_rdata <= 32'hb3a01000;
          16'h0dde : blkif.rom_rdata <= 32'h930e0000;
          16'h0ddf : blkif.rom_rdata <= 32'h130e801f;
          16'h0de0 : blkif.rom_rdata <= 32'h6384d001;
          16'h0de1 : blkif.rom_rdata <= 32'h6f10907e;
          16'h0de2 : blkif.rom_rdata <= 32'hb7000080;
          16'h0de3 : blkif.rom_rdata <= 32'h93804000;
          16'h0de4 : blkif.rom_rdata <= 32'h1301901f;
          16'h0de5 : blkif.rom_rdata <= 32'h23a02000;
          16'h0de6 : blkif.rom_rdata <= 32'h13020000;
          16'h0de7 : blkif.rom_rdata <= 32'h9300b000;
          16'h0de8 : blkif.rom_rdata <= 32'h1301d000;
          16'h0de9 : blkif.rom_rdata <= 32'hb3a12000;
          16'h0dea : blkif.rom_rdata <= 32'h13830100;
          16'h0deb : blkif.rom_rdata <= 32'h13021200;
          16'h0dec : blkif.rom_rdata <= 32'h93022000;
          16'h0ded : blkif.rom_rdata <= 32'he31452fe;
          16'h0dee : blkif.rom_rdata <= 32'h930e1000;
          16'h0def : blkif.rom_rdata <= 32'h130e901f;
          16'h0df0 : blkif.rom_rdata <= 32'h6304d301;
          16'h0df1 : blkif.rom_rdata <= 32'h6f10907a;
          16'h0df2 : blkif.rom_rdata <= 32'hb7000080;
          16'h0df3 : blkif.rom_rdata <= 32'h93804000;
          16'h0df4 : blkif.rom_rdata <= 32'h1301a01f;
          16'h0df5 : blkif.rom_rdata <= 32'h23a02000;
          16'h0df6 : blkif.rom_rdata <= 32'h13020000;
          16'h0df7 : blkif.rom_rdata <= 32'h9300e000;
          16'h0df8 : blkif.rom_rdata <= 32'h1301d000;
          16'h0df9 : blkif.rom_rdata <= 32'hb3a12000;
          16'h0dfa : blkif.rom_rdata <= 32'h13000000;
          16'h0dfb : blkif.rom_rdata <= 32'h13830100;
          16'h0dfc : blkif.rom_rdata <= 32'h13021200;
          16'h0dfd : blkif.rom_rdata <= 32'h93022000;
          16'h0dfe : blkif.rom_rdata <= 32'he31252fe;
          16'h0dff : blkif.rom_rdata <= 32'h930e0000;
          16'h0e00 : blkif.rom_rdata <= 32'h130ea01f;
          16'h0e01 : blkif.rom_rdata <= 32'h6304d301;
          16'h0e02 : blkif.rom_rdata <= 32'h6f105076;
          16'h0e03 : blkif.rom_rdata <= 32'hb7000080;
          16'h0e04 : blkif.rom_rdata <= 32'h93804000;
          16'h0e05 : blkif.rom_rdata <= 32'h1301b01f;
          16'h0e06 : blkif.rom_rdata <= 32'h23a02000;
          16'h0e07 : blkif.rom_rdata <= 32'h13020000;
          16'h0e08 : blkif.rom_rdata <= 32'h9300c000;
          16'h0e09 : blkif.rom_rdata <= 32'h1301d000;
          16'h0e0a : blkif.rom_rdata <= 32'hb3a12000;
          16'h0e0b : blkif.rom_rdata <= 32'h13000000;
          16'h0e0c : blkif.rom_rdata <= 32'h13000000;
          16'h0e0d : blkif.rom_rdata <= 32'h13830100;
          16'h0e0e : blkif.rom_rdata <= 32'h13021200;
          16'h0e0f : blkif.rom_rdata <= 32'h93022000;
          16'h0e10 : blkif.rom_rdata <= 32'he31052fe;
          16'h0e11 : blkif.rom_rdata <= 32'h930e1000;
          16'h0e12 : blkif.rom_rdata <= 32'h130eb01f;
          16'h0e13 : blkif.rom_rdata <= 32'h6304d301;
          16'h0e14 : blkif.rom_rdata <= 32'h6f10d071;
          16'h0e15 : blkif.rom_rdata <= 32'hb7000080;
          16'h0e16 : blkif.rom_rdata <= 32'h93804000;
          16'h0e17 : blkif.rom_rdata <= 32'h1301c01f;
          16'h0e18 : blkif.rom_rdata <= 32'h23a02000;
          16'h0e19 : blkif.rom_rdata <= 32'h13020000;
          16'h0e1a : blkif.rom_rdata <= 32'h9300e000;
          16'h0e1b : blkif.rom_rdata <= 32'h1301d000;
          16'h0e1c : blkif.rom_rdata <= 32'hb3a12000;
          16'h0e1d : blkif.rom_rdata <= 32'h13021200;
          16'h0e1e : blkif.rom_rdata <= 32'h93022000;
          16'h0e1f : blkif.rom_rdata <= 32'he31652fe;
          16'h0e20 : blkif.rom_rdata <= 32'h930e0000;
          16'h0e21 : blkif.rom_rdata <= 32'h130ec01f;
          16'h0e22 : blkif.rom_rdata <= 32'h6384d101;
          16'h0e23 : blkif.rom_rdata <= 32'h6f10106e;
          16'h0e24 : blkif.rom_rdata <= 32'hb7000080;
          16'h0e25 : blkif.rom_rdata <= 32'h93804000;
          16'h0e26 : blkif.rom_rdata <= 32'h1301f01f;
          16'h0e27 : blkif.rom_rdata <= 32'h23a02000;
          16'h0e28 : blkif.rom_rdata <= 32'h13020000;
          16'h0e29 : blkif.rom_rdata <= 32'h9300a000;
          16'h0e2a : blkif.rom_rdata <= 32'h13000000;
          16'h0e2b : blkif.rom_rdata <= 32'h1301d000;
          16'h0e2c : blkif.rom_rdata <= 32'hb3a12000;
          16'h0e2d : blkif.rom_rdata <= 32'h13021200;
          16'h0e2e : blkif.rom_rdata <= 32'h93022000;
          16'h0e2f : blkif.rom_rdata <= 32'he31452fe;
          16'h0e30 : blkif.rom_rdata <= 32'h930e1000;
          16'h0e31 : blkif.rom_rdata <= 32'h130ef01f;
          16'h0e32 : blkif.rom_rdata <= 32'h6384d101;
          16'h0e33 : blkif.rom_rdata <= 32'h6f10106a;
          16'h0e34 : blkif.rom_rdata <= 32'hb7000080;
          16'h0e35 : blkif.rom_rdata <= 32'h93804000;
          16'h0e36 : blkif.rom_rdata <= 32'h13018020;
          16'h0e37 : blkif.rom_rdata <= 32'h23a02000;
          16'h0e38 : blkif.rom_rdata <= 32'h9300f0ff;
          16'h0e39 : blkif.rom_rdata <= 32'h33211000;
          16'h0e3a : blkif.rom_rdata <= 32'h930e0000;
          16'h0e3b : blkif.rom_rdata <= 32'h130e8020;
          16'h0e3c : blkif.rom_rdata <= 32'h6304d101;
          16'h0e3d : blkif.rom_rdata <= 32'h6f109067;
          16'h0e3e : blkif.rom_rdata <= 32'hb7000080;
          16'h0e3f : blkif.rom_rdata <= 32'h93804000;
          16'h0e40 : blkif.rom_rdata <= 32'h13019020;
          16'h0e41 : blkif.rom_rdata <= 32'h23a02000;
          16'h0e42 : blkif.rom_rdata <= 32'h9300f0ff;
          16'h0e43 : blkif.rom_rdata <= 32'h33a10000;
          16'h0e44 : blkif.rom_rdata <= 32'h930e1000;
          16'h0e45 : blkif.rom_rdata <= 32'h130e9020;
          16'h0e46 : blkif.rom_rdata <= 32'h6304d101;
          16'h0e47 : blkif.rom_rdata <= 32'h6f101065;
          16'h0e48 : blkif.rom_rdata <= 32'hb7000080;
          16'h0e49 : blkif.rom_rdata <= 32'h93804000;
          16'h0e4a : blkif.rom_rdata <= 32'h1301a020;
          16'h0e4b : blkif.rom_rdata <= 32'h23a02000;
          16'h0e4c : blkif.rom_rdata <= 32'hb3200000;
          16'h0e4d : blkif.rom_rdata <= 32'h930e0000;
          16'h0e4e : blkif.rom_rdata <= 32'h130ea020;
          16'h0e4f : blkif.rom_rdata <= 32'h6384d001;
          16'h0e50 : blkif.rom_rdata <= 32'h6f10d062;
          16'h0e51 : blkif.rom_rdata <= 32'hb7000080;
          16'h0e52 : blkif.rom_rdata <= 32'h93804000;
          16'h0e53 : blkif.rom_rdata <= 32'h1301b020;
          16'h0e54 : blkif.rom_rdata <= 32'h23a02000;
          16'h0e55 : blkif.rom_rdata <= 32'h93000001;
          16'h0e56 : blkif.rom_rdata <= 32'h1301e001;
          16'h0e57 : blkif.rom_rdata <= 32'h33a02000;
          16'h0e58 : blkif.rom_rdata <= 32'h930e0000;
          16'h0e59 : blkif.rom_rdata <= 32'h130eb020;
          16'h0e5a : blkif.rom_rdata <= 32'h6304d001;
          16'h0e5b : blkif.rom_rdata <= 32'h6f101060;
          16'h0e5c : blkif.rom_rdata <= 32'hb7000080;
          16'h0e5d : blkif.rom_rdata <= 32'h93804000;
          16'h0e5e : blkif.rom_rdata <= 32'h1301c020;
          16'h0e5f : blkif.rom_rdata <= 32'h23a02000;
          16'h0e60 : blkif.rom_rdata <= 32'h93000000;
          16'h0e61 : blkif.rom_rdata <= 32'h93a10000;
          16'h0e62 : blkif.rom_rdata <= 32'h930e0000;
          16'h0e63 : blkif.rom_rdata <= 32'h130ec020;
          16'h0e64 : blkif.rom_rdata <= 32'h6384d101;
          16'h0e65 : blkif.rom_rdata <= 32'h6f10905d;
          16'h0e66 : blkif.rom_rdata <= 32'hb7000080;
          16'h0e67 : blkif.rom_rdata <= 32'h93804000;
          16'h0e68 : blkif.rom_rdata <= 32'h1301e020;
          16'h0e69 : blkif.rom_rdata <= 32'h23a02000;
          16'h0e6a : blkif.rom_rdata <= 32'h93003000;
          16'h0e6b : blkif.rom_rdata <= 32'h93a17000;
          16'h0e6c : blkif.rom_rdata <= 32'h930e1000;
          16'h0e6d : blkif.rom_rdata <= 32'h130ee020;
          16'h0e6e : blkif.rom_rdata <= 32'h6384d101;
          16'h0e6f : blkif.rom_rdata <= 32'h6f10105b;
          16'h0e70 : blkif.rom_rdata <= 32'hb7000080;
          16'h0e71 : blkif.rom_rdata <= 32'h93804000;
          16'h0e72 : blkif.rom_rdata <= 32'h13014021;
          16'h0e73 : blkif.rom_rdata <= 32'h23a02000;
          16'h0e74 : blkif.rom_rdata <= 32'hb7000080;
          16'h0e75 : blkif.rom_rdata <= 32'h9380f0ff;
          16'h0e76 : blkif.rom_rdata <= 32'h93a10000;
          16'h0e77 : blkif.rom_rdata <= 32'h930e0000;
          16'h0e78 : blkif.rom_rdata <= 32'h130e4021;
          16'h0e79 : blkif.rom_rdata <= 32'h6384d101;
          16'h0e7a : blkif.rom_rdata <= 32'h6f105058;
          16'h0e7b : blkif.rom_rdata <= 32'hb7000080;
          16'h0e7c : blkif.rom_rdata <= 32'h93804000;
          16'h0e7d : blkif.rom_rdata <= 32'h13015021;
          16'h0e7e : blkif.rom_rdata <= 32'h23a02000;
          16'h0e7f : blkif.rom_rdata <= 32'hb7000080;
          16'h0e80 : blkif.rom_rdata <= 32'h9380f0ff;
          16'h0e81 : blkif.rom_rdata <= 32'h93a1f07f;
          16'h0e82 : blkif.rom_rdata <= 32'h930e0000;
          16'h0e83 : blkif.rom_rdata <= 32'h130e5021;
          16'h0e84 : blkif.rom_rdata <= 32'h6384d101;
          16'h0e85 : blkif.rom_rdata <= 32'h6f109055;
          16'h0e86 : blkif.rom_rdata <= 32'hb7000080;
          16'h0e87 : blkif.rom_rdata <= 32'h93804000;
          16'h0e88 : blkif.rom_rdata <= 32'h13016021;
          16'h0e89 : blkif.rom_rdata <= 32'h23a02000;
          16'h0e8a : blkif.rom_rdata <= 32'hb7000080;
          16'h0e8b : blkif.rom_rdata <= 32'h93a1f07f;
          16'h0e8c : blkif.rom_rdata <= 32'h930e1000;
          16'h0e8d : blkif.rom_rdata <= 32'h130e6021;
          16'h0e8e : blkif.rom_rdata <= 32'h6384d101;
          16'h0e8f : blkif.rom_rdata <= 32'h6f101053;
          16'h0e90 : blkif.rom_rdata <= 32'hb7000080;
          16'h0e91 : blkif.rom_rdata <= 32'h93804000;
          16'h0e92 : blkif.rom_rdata <= 32'h13017021;
          16'h0e93 : blkif.rom_rdata <= 32'h23a02000;
          16'h0e94 : blkif.rom_rdata <= 32'hb7000080;
          16'h0e95 : blkif.rom_rdata <= 32'h9380f0ff;
          16'h0e96 : blkif.rom_rdata <= 32'h93a10080;
          16'h0e97 : blkif.rom_rdata <= 32'h930e0000;
          16'h0e98 : blkif.rom_rdata <= 32'h130e7021;
          16'h0e99 : blkif.rom_rdata <= 32'h6384d101;
          16'h0e9a : blkif.rom_rdata <= 32'h6f105050;
          16'h0e9b : blkif.rom_rdata <= 32'hb7000080;
          16'h0e9c : blkif.rom_rdata <= 32'h93804000;
          16'h0e9d : blkif.rom_rdata <= 32'h13019021;
          16'h0e9e : blkif.rom_rdata <= 32'h23a02000;
          16'h0e9f : blkif.rom_rdata <= 32'h9300f0ff;
          16'h0ea0 : blkif.rom_rdata <= 32'h93a11000;
          16'h0ea1 : blkif.rom_rdata <= 32'h930e1000;
          16'h0ea2 : blkif.rom_rdata <= 32'h130e9021;
          16'h0ea3 : blkif.rom_rdata <= 32'h6384d101;
          16'h0ea4 : blkif.rom_rdata <= 32'h6f10d04d;
          16'h0ea5 : blkif.rom_rdata <= 32'hb7000080;
          16'h0ea6 : blkif.rom_rdata <= 32'h93804000;
          16'h0ea7 : blkif.rom_rdata <= 32'h1301a021;
          16'h0ea8 : blkif.rom_rdata <= 32'h23a02000;
          16'h0ea9 : blkif.rom_rdata <= 32'h9300f0ff;
          16'h0eaa : blkif.rom_rdata <= 32'h93a1f0ff;
          16'h0eab : blkif.rom_rdata <= 32'h930e0000;
          16'h0eac : blkif.rom_rdata <= 32'h130ea021;
          16'h0ead : blkif.rom_rdata <= 32'h6384d101;
          16'h0eae : blkif.rom_rdata <= 32'h6f10504b;
          16'h0eaf : blkif.rom_rdata <= 32'hb7000080;
          16'h0eb0 : blkif.rom_rdata <= 32'h93804000;
          16'h0eb1 : blkif.rom_rdata <= 32'h1301b021;
          16'h0eb2 : blkif.rom_rdata <= 32'h23a02000;
          16'h0eb3 : blkif.rom_rdata <= 32'h9300b000;
          16'h0eb4 : blkif.rom_rdata <= 32'h93b0d000;
          16'h0eb5 : blkif.rom_rdata <= 32'h930e1000;
          16'h0eb6 : blkif.rom_rdata <= 32'h130eb021;
          16'h0eb7 : blkif.rom_rdata <= 32'h6384d001;
          16'h0eb8 : blkif.rom_rdata <= 32'h6f10d048;
          16'h0eb9 : blkif.rom_rdata <= 32'hb7000080;
          16'h0eba : blkif.rom_rdata <= 32'h93804000;
          16'h0ebb : blkif.rom_rdata <= 32'h1301c021;
          16'h0ebc : blkif.rom_rdata <= 32'h23a02000;
          16'h0ebd : blkif.rom_rdata <= 32'h13020000;
          16'h0ebe : blkif.rom_rdata <= 32'h9300f000;
          16'h0ebf : blkif.rom_rdata <= 32'h93a1a000;
          16'h0ec0 : blkif.rom_rdata <= 32'h13830100;
          16'h0ec1 : blkif.rom_rdata <= 32'h13021200;
          16'h0ec2 : blkif.rom_rdata <= 32'h93022000;
          16'h0ec3 : blkif.rom_rdata <= 32'he31652fe;
          16'h0ec4 : blkif.rom_rdata <= 32'h930e0000;
          16'h0ec5 : blkif.rom_rdata <= 32'h130ec021;
          16'h0ec6 : blkif.rom_rdata <= 32'h6304d301;
          16'h0ec7 : blkif.rom_rdata <= 32'h6f101045;
          16'h0ec8 : blkif.rom_rdata <= 32'hb7000080;
          16'h0ec9 : blkif.rom_rdata <= 32'h93804000;
          16'h0eca : blkif.rom_rdata <= 32'h1301d021;
          16'h0ecb : blkif.rom_rdata <= 32'h23a02000;
          16'h0ecc : blkif.rom_rdata <= 32'h13020000;
          16'h0ecd : blkif.rom_rdata <= 32'h9300a000;
          16'h0ece : blkif.rom_rdata <= 32'h93a10001;
          16'h0ecf : blkif.rom_rdata <= 32'h13000000;
          16'h0ed0 : blkif.rom_rdata <= 32'h13830100;
          16'h0ed1 : blkif.rom_rdata <= 32'h13021200;
          16'h0ed2 : blkif.rom_rdata <= 32'h93022000;
          16'h0ed3 : blkif.rom_rdata <= 32'he31452fe;
          16'h0ed4 : blkif.rom_rdata <= 32'h930e1000;
          16'h0ed5 : blkif.rom_rdata <= 32'h130ed021;
          16'h0ed6 : blkif.rom_rdata <= 32'h6304d301;
          16'h0ed7 : blkif.rom_rdata <= 32'h6f101041;
          16'h0ed8 : blkif.rom_rdata <= 32'hb7000080;
          16'h0ed9 : blkif.rom_rdata <= 32'h93804000;
          16'h0eda : blkif.rom_rdata <= 32'h1301f021;
          16'h0edb : blkif.rom_rdata <= 32'h23a02000;
          16'h0edc : blkif.rom_rdata <= 32'h13020000;
          16'h0edd : blkif.rom_rdata <= 32'h9300b000;
          16'h0ede : blkif.rom_rdata <= 32'h93a1f000;
          16'h0edf : blkif.rom_rdata <= 32'h13021200;
          16'h0ee0 : blkif.rom_rdata <= 32'h93022000;
          16'h0ee1 : blkif.rom_rdata <= 32'he31852fe;
          16'h0ee2 : blkif.rom_rdata <= 32'h930e1000;
          16'h0ee3 : blkif.rom_rdata <= 32'h130ef021;
          16'h0ee4 : blkif.rom_rdata <= 32'h6384d101;
          16'h0ee5 : blkif.rom_rdata <= 32'h6f10903d;
          16'h0ee6 : blkif.rom_rdata <= 32'hb7000080;
          16'h0ee7 : blkif.rom_rdata <= 32'h93804000;
          16'h0ee8 : blkif.rom_rdata <= 32'h13011022;
          16'h0ee9 : blkif.rom_rdata <= 32'h23a02000;
          16'h0eea : blkif.rom_rdata <= 32'h13020000;
          16'h0eeb : blkif.rom_rdata <= 32'h9300c000;
          16'h0eec : blkif.rom_rdata <= 32'h13000000;
          16'h0eed : blkif.rom_rdata <= 32'h13000000;
          16'h0eee : blkif.rom_rdata <= 32'h93a1e000;
          16'h0eef : blkif.rom_rdata <= 32'h13021200;
          16'h0ef0 : blkif.rom_rdata <= 32'h93022000;
          16'h0ef1 : blkif.rom_rdata <= 32'he31452fe;
          16'h0ef2 : blkif.rom_rdata <= 32'h930e1000;
          16'h0ef3 : blkif.rom_rdata <= 32'h130e1022;
          16'h0ef4 : blkif.rom_rdata <= 32'h6384d101;
          16'h0ef5 : blkif.rom_rdata <= 32'h6f109039;
          16'h0ef6 : blkif.rom_rdata <= 32'hb7000080;
          16'h0ef7 : blkif.rom_rdata <= 32'h93804000;
          16'h0ef8 : blkif.rom_rdata <= 32'h13012022;
          16'h0ef9 : blkif.rom_rdata <= 32'h23a02000;
          16'h0efa : blkif.rom_rdata <= 32'h9320f0ff;
          16'h0efb : blkif.rom_rdata <= 32'h930e0000;
          16'h0efc : blkif.rom_rdata <= 32'h130e2022;
          16'h0efd : blkif.rom_rdata <= 32'h6384d001;
          16'h0efe : blkif.rom_rdata <= 32'h6f105037;
          16'h0eff : blkif.rom_rdata <= 32'hb7000080;
          16'h0f00 : blkif.rom_rdata <= 32'h93804000;
          16'h0f01 : blkif.rom_rdata <= 32'h13013022;
          16'h0f02 : blkif.rom_rdata <= 32'h23a02000;
          16'h0f03 : blkif.rom_rdata <= 32'hb700ff00;
          16'h0f04 : blkif.rom_rdata <= 32'h9380f00f;
          16'h0f05 : blkif.rom_rdata <= 32'h13a0f0ff;
          16'h0f06 : blkif.rom_rdata <= 32'h930e0000;
          16'h0f07 : blkif.rom_rdata <= 32'h130e3022;
          16'h0f08 : blkif.rom_rdata <= 32'h6304d001;
          16'h0f09 : blkif.rom_rdata <= 32'h6f109034;
          16'h0f0a : blkif.rom_rdata <= 32'hb7000080;
          16'h0f0b : blkif.rom_rdata <= 32'h93804000;
          16'h0f0c : blkif.rom_rdata <= 32'h13014022;
          16'h0f0d : blkif.rom_rdata <= 32'h23a02000;
          16'h0f0e : blkif.rom_rdata <= 32'hb7000080;
          16'h0f0f : blkif.rom_rdata <= 32'h13010000;
          16'h0f10 : blkif.rom_rdata <= 32'hb3d12040;
          16'h0f11 : blkif.rom_rdata <= 32'hb70e0080;
          16'h0f12 : blkif.rom_rdata <= 32'h130e4022;
          16'h0f13 : blkif.rom_rdata <= 32'h6384d101;
          16'h0f14 : blkif.rom_rdata <= 32'h6f10d031;
          16'h0f15 : blkif.rom_rdata <= 32'hb7000080;
          16'h0f16 : blkif.rom_rdata <= 32'h93804000;
          16'h0f17 : blkif.rom_rdata <= 32'h13015022;
          16'h0f18 : blkif.rom_rdata <= 32'h23a02000;
          16'h0f19 : blkif.rom_rdata <= 32'hb7000080;
          16'h0f1a : blkif.rom_rdata <= 32'h13011000;
          16'h0f1b : blkif.rom_rdata <= 32'hb3d12040;
          16'h0f1c : blkif.rom_rdata <= 32'hb70e00c0;
          16'h0f1d : blkif.rom_rdata <= 32'h130e5022;
          16'h0f1e : blkif.rom_rdata <= 32'h6384d101;
          16'h0f1f : blkif.rom_rdata <= 32'h6f10102f;
          16'h0f20 : blkif.rom_rdata <= 32'hb7000080;
          16'h0f21 : blkif.rom_rdata <= 32'h93804000;
          16'h0f22 : blkif.rom_rdata <= 32'h1301a022;
          16'h0f23 : blkif.rom_rdata <= 32'h23a02000;
          16'h0f24 : blkif.rom_rdata <= 32'hb7000080;
          16'h0f25 : blkif.rom_rdata <= 32'h9380f0ff;
          16'h0f26 : blkif.rom_rdata <= 32'h13011000;
          16'h0f27 : blkif.rom_rdata <= 32'hb3d12040;
          16'h0f28 : blkif.rom_rdata <= 32'hb70e0040;
          16'h0f29 : blkif.rom_rdata <= 32'h938efeff;
          16'h0f2a : blkif.rom_rdata <= 32'h130ea022;
          16'h0f2b : blkif.rom_rdata <= 32'h6384d101;
          16'h0f2c : blkif.rom_rdata <= 32'h6f10d02b;
          16'h0f2d : blkif.rom_rdata <= 32'hb7000080;
          16'h0f2e : blkif.rom_rdata <= 32'h93804000;
          16'h0f2f : blkif.rom_rdata <= 32'h1301f022;
          16'h0f30 : blkif.rom_rdata <= 32'h23a02000;
          16'h0f31 : blkif.rom_rdata <= 32'hb7808181;
          16'h0f32 : blkif.rom_rdata <= 32'h93801018;
          16'h0f33 : blkif.rom_rdata <= 32'h13011000;
          16'h0f34 : blkif.rom_rdata <= 32'hb3d12040;
          16'h0f35 : blkif.rom_rdata <= 32'hb7cec0c0;
          16'h0f36 : blkif.rom_rdata <= 32'h938e0e0c;
          16'h0f37 : blkif.rom_rdata <= 32'h130ef022;
          16'h0f38 : blkif.rom_rdata <= 32'h6384d101;
          16'h0f39 : blkif.rom_rdata <= 32'h6f109028;
          16'h0f3a : blkif.rom_rdata <= 32'hb7000080;
          16'h0f3b : blkif.rom_rdata <= 32'h93804000;
          16'h0f3c : blkif.rom_rdata <= 32'h13013023;
          16'h0f3d : blkif.rom_rdata <= 32'h23a02000;
          16'h0f3e : blkif.rom_rdata <= 32'hb7808181;
          16'h0f3f : blkif.rom_rdata <= 32'h93801018;
          16'h0f40 : blkif.rom_rdata <= 32'h130100fc;
          16'h0f41 : blkif.rom_rdata <= 32'hb3d12040;
          16'h0f42 : blkif.rom_rdata <= 32'hb78e8181;
          16'h0f43 : blkif.rom_rdata <= 32'h938e1e18;
          16'h0f44 : blkif.rom_rdata <= 32'h130e3023;
          16'h0f45 : blkif.rom_rdata <= 32'h6384d101;
          16'h0f46 : blkif.rom_rdata <= 32'h6f105025;
          16'h0f47 : blkif.rom_rdata <= 32'hb7000080;
          16'h0f48 : blkif.rom_rdata <= 32'h93804000;
          16'h0f49 : blkif.rom_rdata <= 32'h13016023;
          16'h0f4a : blkif.rom_rdata <= 32'h23a02000;
          16'h0f4b : blkif.rom_rdata <= 32'hb7808181;
          16'h0f4c : blkif.rom_rdata <= 32'h93801018;
          16'h0f4d : blkif.rom_rdata <= 32'h1301e0fc;
          16'h0f4e : blkif.rom_rdata <= 32'hb3d12040;
          16'h0f4f : blkif.rom_rdata <= 32'hb70efeff;
          16'h0f50 : blkif.rom_rdata <= 32'h938e6e60;
          16'h0f51 : blkif.rom_rdata <= 32'h130e6023;
          16'h0f52 : blkif.rom_rdata <= 32'h6384d101;
          16'h0f53 : blkif.rom_rdata <= 32'h6f101022;
          16'h0f54 : blkif.rom_rdata <= 32'hb7000080;
          16'h0f55 : blkif.rom_rdata <= 32'h93804000;
          16'h0f56 : blkif.rom_rdata <= 32'h13017023;
          16'h0f57 : blkif.rom_rdata <= 32'h23a02000;
          16'h0f58 : blkif.rom_rdata <= 32'hb7808181;
          16'h0f59 : blkif.rom_rdata <= 32'h93801018;
          16'h0f5a : blkif.rom_rdata <= 32'h1301f0ff;
          16'h0f5b : blkif.rom_rdata <= 32'hb3d12040;
          16'h0f5c : blkif.rom_rdata <= 32'h930ef0ff;
          16'h0f5d : blkif.rom_rdata <= 32'h130e7023;
          16'h0f5e : blkif.rom_rdata <= 32'h6384d101;
          16'h0f5f : blkif.rom_rdata <= 32'h6f10101f;
          16'h0f60 : blkif.rom_rdata <= 32'hb7000080;
          16'h0f61 : blkif.rom_rdata <= 32'h93804000;
          16'h0f62 : blkif.rom_rdata <= 32'h13018023;
          16'h0f63 : blkif.rom_rdata <= 32'h23a02000;
          16'h0f64 : blkif.rom_rdata <= 32'hb7000080;
          16'h0f65 : blkif.rom_rdata <= 32'h13017000;
          16'h0f66 : blkif.rom_rdata <= 32'hb3d02040;
          16'h0f67 : blkif.rom_rdata <= 32'hb70e00ff;
          16'h0f68 : blkif.rom_rdata <= 32'h130e8023;
          16'h0f69 : blkif.rom_rdata <= 32'h6384d001;
          16'h0f6a : blkif.rom_rdata <= 32'h6f10501c;
          16'h0f6b : blkif.rom_rdata <= 32'hb7000080;
          16'h0f6c : blkif.rom_rdata <= 32'h93804000;
          16'h0f6d : blkif.rom_rdata <= 32'h13019023;
          16'h0f6e : blkif.rom_rdata <= 32'h23a02000;
          16'h0f6f : blkif.rom_rdata <= 32'hb7000080;
          16'h0f70 : blkif.rom_rdata <= 32'h1301e000;
          16'h0f71 : blkif.rom_rdata <= 32'h33d12040;
          16'h0f72 : blkif.rom_rdata <= 32'hb70efeff;
          16'h0f73 : blkif.rom_rdata <= 32'h130e9023;
          16'h0f74 : blkif.rom_rdata <= 32'h6304d101;
          16'h0f75 : blkif.rom_rdata <= 32'h6f109019;
          16'h0f76 : blkif.rom_rdata <= 32'hb7000080;
          16'h0f77 : blkif.rom_rdata <= 32'h93804000;
          16'h0f78 : blkif.rom_rdata <= 32'h1301a023;
          16'h0f79 : blkif.rom_rdata <= 32'h23a02000;
          16'h0f7a : blkif.rom_rdata <= 32'h93007000;
          16'h0f7b : blkif.rom_rdata <= 32'hb3d01040;
          16'h0f7c : blkif.rom_rdata <= 32'h930e0000;
          16'h0f7d : blkif.rom_rdata <= 32'h130ea023;
          16'h0f7e : blkif.rom_rdata <= 32'h6384d001;
          16'h0f7f : blkif.rom_rdata <= 32'h6f101017;
          16'h0f80 : blkif.rom_rdata <= 32'hb7000080;
          16'h0f81 : blkif.rom_rdata <= 32'h93804000;
          16'h0f82 : blkif.rom_rdata <= 32'h1301b023;
          16'h0f83 : blkif.rom_rdata <= 32'h23a02000;
          16'h0f84 : blkif.rom_rdata <= 32'h13020000;
          16'h0f85 : blkif.rom_rdata <= 32'hb7000080;
          16'h0f86 : blkif.rom_rdata <= 32'h13017000;
          16'h0f87 : blkif.rom_rdata <= 32'hb3d12040;
          16'h0f88 : blkif.rom_rdata <= 32'h13830100;
          16'h0f89 : blkif.rom_rdata <= 32'h13021200;
          16'h0f8a : blkif.rom_rdata <= 32'h93022000;
          16'h0f8b : blkif.rom_rdata <= 32'he31452fe;
          16'h0f8c : blkif.rom_rdata <= 32'hb70e00ff;
          16'h0f8d : blkif.rom_rdata <= 32'h130eb023;
          16'h0f8e : blkif.rom_rdata <= 32'h6304d301;
          16'h0f8f : blkif.rom_rdata <= 32'h6f101013;
          16'h0f90 : blkif.rom_rdata <= 32'hb7000080;
          16'h0f91 : blkif.rom_rdata <= 32'h93804000;
          16'h0f92 : blkif.rom_rdata <= 32'h1301c023;
          16'h0f93 : blkif.rom_rdata <= 32'h23a02000;
          16'h0f94 : blkif.rom_rdata <= 32'h13020000;
          16'h0f95 : blkif.rom_rdata <= 32'hb7000080;
          16'h0f96 : blkif.rom_rdata <= 32'h1301e000;
          16'h0f97 : blkif.rom_rdata <= 32'hb3d12040;
          16'h0f98 : blkif.rom_rdata <= 32'h13000000;
          16'h0f99 : blkif.rom_rdata <= 32'h13830100;
          16'h0f9a : blkif.rom_rdata <= 32'h13021200;
          16'h0f9b : blkif.rom_rdata <= 32'h93022000;
          16'h0f9c : blkif.rom_rdata <= 32'he31252fe;
          16'h0f9d : blkif.rom_rdata <= 32'hb70efeff;
          16'h0f9e : blkif.rom_rdata <= 32'h130ec023;
          16'h0f9f : blkif.rom_rdata <= 32'h6304d301;
          16'h0fa0 : blkif.rom_rdata <= 32'h6f10d00e;
          16'h0fa1 : blkif.rom_rdata <= 32'hb7000080;
          16'h0fa2 : blkif.rom_rdata <= 32'h93804000;
          16'h0fa3 : blkif.rom_rdata <= 32'h13014024;
          16'h0fa4 : blkif.rom_rdata <= 32'h23a02000;
          16'h0fa5 : blkif.rom_rdata <= 32'h13020000;
          16'h0fa6 : blkif.rom_rdata <= 32'h13017000;
          16'h0fa7 : blkif.rom_rdata <= 32'hb7000080;
          16'h0fa8 : blkif.rom_rdata <= 32'hb3d12040;
          16'h0fa9 : blkif.rom_rdata <= 32'h13021200;
          16'h0faa : blkif.rom_rdata <= 32'h93022000;
          16'h0fab : blkif.rom_rdata <= 32'he31652fe;
          16'h0fac : blkif.rom_rdata <= 32'hb70e00ff;
          16'h0fad : blkif.rom_rdata <= 32'h130e4024;
          16'h0fae : blkif.rom_rdata <= 32'h6384d101;
          16'h0faf : blkif.rom_rdata <= 32'h6f10100b;
          16'h0fb0 : blkif.rom_rdata <= 32'hb7000080;
          16'h0fb1 : blkif.rom_rdata <= 32'h93804000;
          16'h0fb2 : blkif.rom_rdata <= 32'h13019024;
          16'h0fb3 : blkif.rom_rdata <= 32'h23a02000;
          16'h0fb4 : blkif.rom_rdata <= 32'h13020000;
          16'h0fb5 : blkif.rom_rdata <= 32'h1301f001;
          16'h0fb6 : blkif.rom_rdata <= 32'h13000000;
          16'h0fb7 : blkif.rom_rdata <= 32'h13000000;
          16'h0fb8 : blkif.rom_rdata <= 32'hb7000080;
          16'h0fb9 : blkif.rom_rdata <= 32'hb3d12040;
          16'h0fba : blkif.rom_rdata <= 32'h13021200;
          16'h0fbb : blkif.rom_rdata <= 32'h93022000;
          16'h0fbc : blkif.rom_rdata <= 32'he31252fe;
          16'h0fbd : blkif.rom_rdata <= 32'h930ef0ff;
          16'h0fbe : blkif.rom_rdata <= 32'h130e9024;
          16'h0fbf : blkif.rom_rdata <= 32'h6384d101;
          16'h0fc0 : blkif.rom_rdata <= 32'h6f10d006;
          16'h0fc1 : blkif.rom_rdata <= 32'hb7000080;
          16'h0fc2 : blkif.rom_rdata <= 32'h93804000;
          16'h0fc3 : blkif.rom_rdata <= 32'h1301a024;
          16'h0fc4 : blkif.rom_rdata <= 32'h23a02000;
          16'h0fc5 : blkif.rom_rdata <= 32'h9300f000;
          16'h0fc6 : blkif.rom_rdata <= 32'h33511040;
          16'h0fc7 : blkif.rom_rdata <= 32'h930e0000;
          16'h0fc8 : blkif.rom_rdata <= 32'h130ea024;
          16'h0fc9 : blkif.rom_rdata <= 32'h6304d101;
          16'h0fca : blkif.rom_rdata <= 32'h6f105004;
          16'h0fcb : blkif.rom_rdata <= 32'hb7000080;
          16'h0fcc : blkif.rom_rdata <= 32'h93804000;
          16'h0fcd : blkif.rom_rdata <= 32'h1301b024;
          16'h0fce : blkif.rom_rdata <= 32'h23a02000;
          16'h0fcf : blkif.rom_rdata <= 32'h93000002;
          16'h0fd0 : blkif.rom_rdata <= 32'h33d10040;
          16'h0fd1 : blkif.rom_rdata <= 32'h930e0002;
          16'h0fd2 : blkif.rom_rdata <= 32'h130eb024;
          16'h0fd3 : blkif.rom_rdata <= 32'h6304d101;
          16'h0fd4 : blkif.rom_rdata <= 32'h6f10d001;
          16'h0fd5 : blkif.rom_rdata <= 32'hb7000080;
          16'h0fd6 : blkif.rom_rdata <= 32'h93804000;
          16'h0fd7 : blkif.rom_rdata <= 32'h1301c024;
          16'h0fd8 : blkif.rom_rdata <= 32'h23a02000;
          16'h0fd9 : blkif.rom_rdata <= 32'hb3500040;
          16'h0fda : blkif.rom_rdata <= 32'h930e0000;
          16'h0fdb : blkif.rom_rdata <= 32'h130ec024;
          16'h0fdc : blkif.rom_rdata <= 32'h6384d001;
          16'h0fdd : blkif.rom_rdata <= 32'h6f10807f;
          16'h0fde : blkif.rom_rdata <= 32'hb7000080;
          16'h0fdf : blkif.rom_rdata <= 32'h93804000;
          16'h0fe0 : blkif.rom_rdata <= 32'h1301d024;
          16'h0fe1 : blkif.rom_rdata <= 32'h23a02000;
          16'h0fe2 : blkif.rom_rdata <= 32'h93000040;
          16'h0fe3 : blkif.rom_rdata <= 32'h37110000;
          16'h0fe4 : blkif.rom_rdata <= 32'h13010180;
          16'h0fe5 : blkif.rom_rdata <= 32'h33d02040;
          16'h0fe6 : blkif.rom_rdata <= 32'h930e0000;
          16'h0fe7 : blkif.rom_rdata <= 32'h130ed024;
          16'h0fe8 : blkif.rom_rdata <= 32'h6304d001;
          16'h0fe9 : blkif.rom_rdata <= 32'h6f10807c;
          16'h0fea : blkif.rom_rdata <= 32'hb7000080;
          16'h0feb : blkif.rom_rdata <= 32'h93804000;
          16'h0fec : blkif.rom_rdata <= 32'h1301e024;
          16'h0fed : blkif.rom_rdata <= 32'h23a02000;
          16'h0fee : blkif.rom_rdata <= 32'h93000000;
          16'h0fef : blkif.rom_rdata <= 32'h93d10040;
          16'h0ff0 : blkif.rom_rdata <= 32'h930e0000;
          16'h0ff1 : blkif.rom_rdata <= 32'h130ee024;
          16'h0ff2 : blkif.rom_rdata <= 32'h6384d101;
          16'h0ff3 : blkif.rom_rdata <= 32'h6f10007a;
          16'h0ff4 : blkif.rom_rdata <= 32'hb7000080;
          16'h0ff5 : blkif.rom_rdata <= 32'h93804000;
          16'h0ff6 : blkif.rom_rdata <= 32'h13015025;
          16'h0ff7 : blkif.rom_rdata <= 32'h23a02000;
          16'h0ff8 : blkif.rom_rdata <= 32'hb7000080;
          16'h0ff9 : blkif.rom_rdata <= 32'h9380f0ff;
          16'h0ffa : blkif.rom_rdata <= 32'h93d17040;
          16'h0ffb : blkif.rom_rdata <= 32'hb70e0001;
          16'h0ffc : blkif.rom_rdata <= 32'h938efeff;
          16'h0ffd : blkif.rom_rdata <= 32'h130e5025;
          16'h0ffe : blkif.rom_rdata <= 32'h6384d101;
          16'h0fff : blkif.rom_rdata <= 32'h6f100077;
          16'h1000 : blkif.rom_rdata <= 32'hb7000080;
          16'h1001 : blkif.rom_rdata <= 32'h93804000;
          16'h1002 : blkif.rom_rdata <= 32'h13017025;
          16'h1003 : blkif.rom_rdata <= 32'h23a02000;
          16'h1004 : blkif.rom_rdata <= 32'hb7000080;
          16'h1005 : blkif.rom_rdata <= 32'h9380f0ff;
          16'h1006 : blkif.rom_rdata <= 32'h93d1f041;
          16'h1007 : blkif.rom_rdata <= 32'h930e0000;
          16'h1008 : blkif.rom_rdata <= 32'h130e7025;
          16'h1009 : blkif.rom_rdata <= 32'h6384d101;
          16'h100a : blkif.rom_rdata <= 32'h6f104074;
          16'h100b : blkif.rom_rdata <= 32'hb7000080;
          16'h100c : blkif.rom_rdata <= 32'h93804000;
          16'h100d : blkif.rom_rdata <= 32'h13018025;
          16'h100e : blkif.rom_rdata <= 32'h23a02000;
          16'h100f : blkif.rom_rdata <= 32'hb7808181;
          16'h1010 : blkif.rom_rdata <= 32'h93801018;
          16'h1011 : blkif.rom_rdata <= 32'h93d10040;
          16'h1012 : blkif.rom_rdata <= 32'hb78e8181;
          16'h1013 : blkif.rom_rdata <= 32'h938e1e18;
          16'h1014 : blkif.rom_rdata <= 32'h130e8025;
          16'h1015 : blkif.rom_rdata <= 32'h6384d101;
          16'h1016 : blkif.rom_rdata <= 32'h6f104071;
          16'h1017 : blkif.rom_rdata <= 32'hb7000080;
          16'h1018 : blkif.rom_rdata <= 32'h93804000;
          16'h1019 : blkif.rom_rdata <= 32'h13019025;
          16'h101a : blkif.rom_rdata <= 32'h23a02000;
          16'h101b : blkif.rom_rdata <= 32'hb7808181;
          16'h101c : blkif.rom_rdata <= 32'h93801018;
          16'h101d : blkif.rom_rdata <= 32'h93d11040;
          16'h101e : blkif.rom_rdata <= 32'hb7cec0c0;
          16'h101f : blkif.rom_rdata <= 32'h938e0e0c;
          16'h1020 : blkif.rom_rdata <= 32'h130e9025;
          16'h1021 : blkif.rom_rdata <= 32'h6384d101;
          16'h1022 : blkif.rom_rdata <= 32'h6f10406e;
          16'h1023 : blkif.rom_rdata <= 32'hb7000080;
          16'h1024 : blkif.rom_rdata <= 32'h93804000;
          16'h1025 : blkif.rom_rdata <= 32'h1301d025;
          16'h1026 : blkif.rom_rdata <= 32'h23a02000;
          16'h1027 : blkif.rom_rdata <= 32'hb7000080;
          16'h1028 : blkif.rom_rdata <= 32'h93d07040;
          16'h1029 : blkif.rom_rdata <= 32'hb70e00ff;
          16'h102a : blkif.rom_rdata <= 32'h130ed025;
          16'h102b : blkif.rom_rdata <= 32'h6384d001;
          16'h102c : blkif.rom_rdata <= 32'h6f10c06b;
          16'h102d : blkif.rom_rdata <= 32'hb7000080;
          16'h102e : blkif.rom_rdata <= 32'h93804000;
          16'h102f : blkif.rom_rdata <= 32'h1301e025;
          16'h1030 : blkif.rom_rdata <= 32'h23a02000;
          16'h1031 : blkif.rom_rdata <= 32'h13020000;
          16'h1032 : blkif.rom_rdata <= 32'hb7000080;
          16'h1033 : blkif.rom_rdata <= 32'h93d17040;
          16'h1034 : blkif.rom_rdata <= 32'h13830100;
          16'h1035 : blkif.rom_rdata <= 32'h13021200;
          16'h1036 : blkif.rom_rdata <= 32'h93022000;
          16'h1037 : blkif.rom_rdata <= 32'he31652fe;
          16'h1038 : blkif.rom_rdata <= 32'hb70e00ff;
          16'h1039 : blkif.rom_rdata <= 32'h130ee025;
          16'h103a : blkif.rom_rdata <= 32'h6304d301;
          16'h103b : blkif.rom_rdata <= 32'h6f100068;
          16'h103c : blkif.rom_rdata <= 32'hb7000080;
          16'h103d : blkif.rom_rdata <= 32'h93804000;
          16'h103e : blkif.rom_rdata <= 32'h13011026;
          16'h103f : blkif.rom_rdata <= 32'h23a02000;
          16'h1040 : blkif.rom_rdata <= 32'h13020000;
          16'h1041 : blkif.rom_rdata <= 32'hb7000080;
          16'h1042 : blkif.rom_rdata <= 32'h93d17040;
          16'h1043 : blkif.rom_rdata <= 32'h13021200;
          16'h1044 : blkif.rom_rdata <= 32'h93022000;
          16'h1045 : blkif.rom_rdata <= 32'he31852fe;
          16'h1046 : blkif.rom_rdata <= 32'hb70e00ff;
          16'h1047 : blkif.rom_rdata <= 32'h130e1026;
          16'h1048 : blkif.rom_rdata <= 32'h6384d101;
          16'h1049 : blkif.rom_rdata <= 32'h6f108064;
          16'h104a : blkif.rom_rdata <= 32'hb7000080;
          16'h104b : blkif.rom_rdata <= 32'h93804000;
          16'h104c : blkif.rom_rdata <= 32'h13012026;
          16'h104d : blkif.rom_rdata <= 32'h23a02000;
          16'h104e : blkif.rom_rdata <= 32'h13020000;
          16'h104f : blkif.rom_rdata <= 32'hb7000080;
          16'h1050 : blkif.rom_rdata <= 32'h13000000;
          16'h1051 : blkif.rom_rdata <= 32'h93d1e040;
          16'h1052 : blkif.rom_rdata <= 32'h13021200;
          16'h1053 : blkif.rom_rdata <= 32'h93022000;
          16'h1054 : blkif.rom_rdata <= 32'he31652fe;
          16'h1055 : blkif.rom_rdata <= 32'hb70efeff;
          16'h1056 : blkif.rom_rdata <= 32'h130e2026;
          16'h1057 : blkif.rom_rdata <= 32'h6384d101;
          16'h1058 : blkif.rom_rdata <= 32'h6f10c060;
          16'h1059 : blkif.rom_rdata <= 32'hb7000080;
          16'h105a : blkif.rom_rdata <= 32'h93804000;
          16'h105b : blkif.rom_rdata <= 32'h13014026;
          16'h105c : blkif.rom_rdata <= 32'h23a02000;
          16'h105d : blkif.rom_rdata <= 32'h9350f041;
          16'h105e : blkif.rom_rdata <= 32'h930e0000;
          16'h105f : blkif.rom_rdata <= 32'h130e4026;
          16'h1060 : blkif.rom_rdata <= 32'h6384d001;
          16'h1061 : blkif.rom_rdata <= 32'h6f10805e;
          16'h1062 : blkif.rom_rdata <= 32'hb7000080;
          16'h1063 : blkif.rom_rdata <= 32'h93804000;
          16'h1064 : blkif.rom_rdata <= 32'h13015026;
          16'h1065 : blkif.rom_rdata <= 32'h23a02000;
          16'h1066 : blkif.rom_rdata <= 32'h93001002;
          16'h1067 : blkif.rom_rdata <= 32'h13d04041;
          16'h1068 : blkif.rom_rdata <= 32'h930e0000;
          16'h1069 : blkif.rom_rdata <= 32'h130e5026;
          16'h106a : blkif.rom_rdata <= 32'h6304d001;
          16'h106b : blkif.rom_rdata <= 32'h6f10005c;
          16'h106c : blkif.rom_rdata <= 32'hb7000080;
          16'h106d : blkif.rom_rdata <= 32'h93804000;
          16'h106e : blkif.rom_rdata <= 32'h13016026;
          16'h106f : blkif.rom_rdata <= 32'h23a02000;
          16'h1070 : blkif.rom_rdata <= 32'hb780ffff;
          16'h1071 : blkif.rom_rdata <= 32'h13010000;
          16'h1072 : blkif.rom_rdata <= 32'hb3d12000;
          16'h1073 : blkif.rom_rdata <= 32'hb78effff;
          16'h1074 : blkif.rom_rdata <= 32'h130e6026;
          16'h1075 : blkif.rom_rdata <= 32'h6384d101;
          16'h1076 : blkif.rom_rdata <= 32'h6f104059;
          16'h1077 : blkif.rom_rdata <= 32'hb7000080;
          16'h1078 : blkif.rom_rdata <= 32'h93804000;
          16'h1079 : blkif.rom_rdata <= 32'h1301b026;
          16'h107a : blkif.rom_rdata <= 32'h23a02000;
          16'h107b : blkif.rom_rdata <= 32'h9300f0ff;
          16'h107c : blkif.rom_rdata <= 32'h13010000;
          16'h107d : blkif.rom_rdata <= 32'hb3d12000;
          16'h107e : blkif.rom_rdata <= 32'h930ef0ff;
          16'h107f : blkif.rom_rdata <= 32'h130eb026;
          16'h1080 : blkif.rom_rdata <= 32'h6384d101;
          16'h1081 : blkif.rom_rdata <= 32'h6f108056;
          16'h1082 : blkif.rom_rdata <= 32'hb7000080;
          16'h1083 : blkif.rom_rdata <= 32'h93804000;
          16'h1084 : blkif.rom_rdata <= 32'h1301f026;
          16'h1085 : blkif.rom_rdata <= 32'h23a02000;
          16'h1086 : blkif.rom_rdata <= 32'h9300f0ff;
          16'h1087 : blkif.rom_rdata <= 32'h1301f001;
          16'h1088 : blkif.rom_rdata <= 32'hb3d12000;
          16'h1089 : blkif.rom_rdata <= 32'h930e1000;
          16'h108a : blkif.rom_rdata <= 32'h130ef026;
          16'h108b : blkif.rom_rdata <= 32'h6384d101;
          16'h108c : blkif.rom_rdata <= 32'h6f10c053;
          16'h108d : blkif.rom_rdata <= 32'hb7000080;
          16'h108e : blkif.rom_rdata <= 32'h93804000;
          16'h108f : blkif.rom_rdata <= 32'h13010027;
          16'h1090 : blkif.rom_rdata <= 32'h23a02000;
          16'h1091 : blkif.rom_rdata <= 32'hb7202121;
          16'h1092 : blkif.rom_rdata <= 32'h93801012;
          16'h1093 : blkif.rom_rdata <= 32'h13010000;
          16'h1094 : blkif.rom_rdata <= 32'hb3d12000;
          16'h1095 : blkif.rom_rdata <= 32'hb72e2121;
          16'h1096 : blkif.rom_rdata <= 32'h938e1e12;
          16'h1097 : blkif.rom_rdata <= 32'h130e0027;
          16'h1098 : blkif.rom_rdata <= 32'h6384d101;
          16'h1099 : blkif.rom_rdata <= 32'h6f108050;
          16'h109a : blkif.rom_rdata <= 32'hb7000080;
          16'h109b : blkif.rom_rdata <= 32'h93804000;
          16'h109c : blkif.rom_rdata <= 32'h13015027;
          16'h109d : blkif.rom_rdata <= 32'h23a02000;
          16'h109e : blkif.rom_rdata <= 32'hb7202121;
          16'h109f : blkif.rom_rdata <= 32'h93801012;
          16'h10a0 : blkif.rom_rdata <= 32'h130100fe;
          16'h10a1 : blkif.rom_rdata <= 32'hb3d12000;
          16'h10a2 : blkif.rom_rdata <= 32'hb72e2121;
          16'h10a3 : blkif.rom_rdata <= 32'h938e1e12;
          16'h10a4 : blkif.rom_rdata <= 32'h130e5027;
          16'h10a5 : blkif.rom_rdata <= 32'h6384d101;
          16'h10a6 : blkif.rom_rdata <= 32'h6f10404d;
          16'h10a7 : blkif.rom_rdata <= 32'hb7000080;
          16'h10a8 : blkif.rom_rdata <= 32'h93804000;
          16'h10a9 : blkif.rom_rdata <= 32'h13016027;
          16'h10aa : blkif.rom_rdata <= 32'h23a02000;
          16'h10ab : blkif.rom_rdata <= 32'hb7202121;
          16'h10ac : blkif.rom_rdata <= 32'h93801012;
          16'h10ad : blkif.rom_rdata <= 32'h130110fe;
          16'h10ae : blkif.rom_rdata <= 32'hb3d12000;
          16'h10af : blkif.rom_rdata <= 32'hb79e9010;
          16'h10b0 : blkif.rom_rdata <= 32'h938e0e09;
          16'h10b1 : blkif.rom_rdata <= 32'h130e6027;
          16'h10b2 : blkif.rom_rdata <= 32'h6384d101;
          16'h10b3 : blkif.rom_rdata <= 32'h6f10004a;
          16'h10b4 : blkif.rom_rdata <= 32'hb7000080;
          16'h10b5 : blkif.rom_rdata <= 32'h93804000;
          16'h10b6 : blkif.rom_rdata <= 32'h13017027;
          16'h10b7 : blkif.rom_rdata <= 32'h23a02000;
          16'h10b8 : blkif.rom_rdata <= 32'hb7202121;
          16'h10b9 : blkif.rom_rdata <= 32'h93801012;
          16'h10ba : blkif.rom_rdata <= 32'h130170fe;
          16'h10bb : blkif.rom_rdata <= 32'hb3d12000;
          16'h10bc : blkif.rom_rdata <= 32'hb74e4200;
          16'h10bd : blkif.rom_rdata <= 32'h938e2e24;
          16'h10be : blkif.rom_rdata <= 32'h130e7027;
          16'h10bf : blkif.rom_rdata <= 32'h6384d101;
          16'h10c0 : blkif.rom_rdata <= 32'h6f10c046;
          16'h10c1 : blkif.rom_rdata <= 32'hb7000080;
          16'h10c2 : blkif.rom_rdata <= 32'h93804000;
          16'h10c3 : blkif.rom_rdata <= 32'h1301a027;
          16'h10c4 : blkif.rom_rdata <= 32'h23a02000;
          16'h10c5 : blkif.rom_rdata <= 32'hb780ffff;
          16'h10c6 : blkif.rom_rdata <= 32'h13011000;
          16'h10c7 : blkif.rom_rdata <= 32'hb3d02000;
          16'h10c8 : blkif.rom_rdata <= 32'hb7ceff7f;
          16'h10c9 : blkif.rom_rdata <= 32'h130ea027;
          16'h10ca : blkif.rom_rdata <= 32'h6384d001;
          16'h10cb : blkif.rom_rdata <= 32'h6f100044;
          16'h10cc : blkif.rom_rdata <= 32'hb7000080;
          16'h10cd : blkif.rom_rdata <= 32'h93804000;
          16'h10ce : blkif.rom_rdata <= 32'h1301b027;
          16'h10cf : blkif.rom_rdata <= 32'h23a02000;
          16'h10d0 : blkif.rom_rdata <= 32'hb780ffff;
          16'h10d1 : blkif.rom_rdata <= 32'h1301e000;
          16'h10d2 : blkif.rom_rdata <= 32'h33d12000;
          16'h10d3 : blkif.rom_rdata <= 32'hb70e0400;
          16'h10d4 : blkif.rom_rdata <= 32'h938eeeff;
          16'h10d5 : blkif.rom_rdata <= 32'h130eb027;
          16'h10d6 : blkif.rom_rdata <= 32'h6304d101;
          16'h10d7 : blkif.rom_rdata <= 32'h6f100041;
          16'h10d8 : blkif.rom_rdata <= 32'hb7000080;
          16'h10d9 : blkif.rom_rdata <= 32'h93804000;
          16'h10da : blkif.rom_rdata <= 32'h1301c027;
          16'h10db : blkif.rom_rdata <= 32'h23a02000;
          16'h10dc : blkif.rom_rdata <= 32'h93007000;
          16'h10dd : blkif.rom_rdata <= 32'hb3d01000;
          16'h10de : blkif.rom_rdata <= 32'h930e0000;
          16'h10df : blkif.rom_rdata <= 32'h130ec027;
          16'h10e0 : blkif.rom_rdata <= 32'h6384d001;
          16'h10e1 : blkif.rom_rdata <= 32'h6f10803e;
          16'h10e2 : blkif.rom_rdata <= 32'hb7000080;
          16'h10e3 : blkif.rom_rdata <= 32'h93804000;
          16'h10e4 : blkif.rom_rdata <= 32'h1301d027;
          16'h10e5 : blkif.rom_rdata <= 32'h23a02000;
          16'h10e6 : blkif.rom_rdata <= 32'h13020000;
          16'h10e7 : blkif.rom_rdata <= 32'hb780ffff;
          16'h10e8 : blkif.rom_rdata <= 32'h13011000;
          16'h10e9 : blkif.rom_rdata <= 32'hb3d12000;
          16'h10ea : blkif.rom_rdata <= 32'h13830100;
          16'h10eb : blkif.rom_rdata <= 32'h13021200;
          16'h10ec : blkif.rom_rdata <= 32'h93022000;
          16'h10ed : blkif.rom_rdata <= 32'he31452fe;
          16'h10ee : blkif.rom_rdata <= 32'hb7ceff7f;
          16'h10ef : blkif.rom_rdata <= 32'h130ed027;
          16'h10f0 : blkif.rom_rdata <= 32'h6304d301;
          16'h10f1 : blkif.rom_rdata <= 32'h6f10803a;
          16'h10f2 : blkif.rom_rdata <= 32'hb7000080;
          16'h10f3 : blkif.rom_rdata <= 32'h93804000;
          16'h10f4 : blkif.rom_rdata <= 32'h13010028;
          16'h10f5 : blkif.rom_rdata <= 32'h23a02000;
          16'h10f6 : blkif.rom_rdata <= 32'h13020000;
          16'h10f7 : blkif.rom_rdata <= 32'hb780ffff;
          16'h10f8 : blkif.rom_rdata <= 32'h13011000;
          16'h10f9 : blkif.rom_rdata <= 32'hb3d12000;
          16'h10fa : blkif.rom_rdata <= 32'h13021200;
          16'h10fb : blkif.rom_rdata <= 32'h93022000;
          16'h10fc : blkif.rom_rdata <= 32'he31652fe;
          16'h10fd : blkif.rom_rdata <= 32'hb7ceff7f;
          16'h10fe : blkif.rom_rdata <= 32'h130e0028;
          16'h10ff : blkif.rom_rdata <= 32'h6384d101;
          16'h1100 : blkif.rom_rdata <= 32'h6f10c036;
          16'h1101 : blkif.rom_rdata <= 32'hb7000080;
          16'h1102 : blkif.rom_rdata <= 32'h93804000;
          16'h1103 : blkif.rom_rdata <= 32'h13016028;
          16'h1104 : blkif.rom_rdata <= 32'h23a02000;
          16'h1105 : blkif.rom_rdata <= 32'h13020000;
          16'h1106 : blkif.rom_rdata <= 32'h13011000;
          16'h1107 : blkif.rom_rdata <= 32'hb780ffff;
          16'h1108 : blkif.rom_rdata <= 32'hb3d12000;
          16'h1109 : blkif.rom_rdata <= 32'h13021200;
          16'h110a : blkif.rom_rdata <= 32'h93022000;
          16'h110b : blkif.rom_rdata <= 32'he31652fe;
          16'h110c : blkif.rom_rdata <= 32'hb7ceff7f;
          16'h110d : blkif.rom_rdata <= 32'h130e6028;
          16'h110e : blkif.rom_rdata <= 32'h6384d101;
          16'h110f : blkif.rom_rdata <= 32'h6f100033;
          16'h1110 : blkif.rom_rdata <= 32'hb7000080;
          16'h1111 : blkif.rom_rdata <= 32'h93804000;
          16'h1112 : blkif.rom_rdata <= 32'h1301b028;
          16'h1113 : blkif.rom_rdata <= 32'h23a02000;
          16'h1114 : blkif.rom_rdata <= 32'h13020000;
          16'h1115 : blkif.rom_rdata <= 32'h1301f000;
          16'h1116 : blkif.rom_rdata <= 32'h13000000;
          16'h1117 : blkif.rom_rdata <= 32'h13000000;
          16'h1118 : blkif.rom_rdata <= 32'hb780ffff;
          16'h1119 : blkif.rom_rdata <= 32'hb3d12000;
          16'h111a : blkif.rom_rdata <= 32'h13021200;
          16'h111b : blkif.rom_rdata <= 32'h93022000;
          16'h111c : blkif.rom_rdata <= 32'he31252fe;
          16'h111d : blkif.rom_rdata <= 32'hb70e0200;
          16'h111e : blkif.rom_rdata <= 32'h938efeff;
          16'h111f : blkif.rom_rdata <= 32'h130eb028;
          16'h1120 : blkif.rom_rdata <= 32'h6384d101;
          16'h1121 : blkif.rom_rdata <= 32'h6f10802e;
          16'h1122 : blkif.rom_rdata <= 32'hb7000080;
          16'h1123 : blkif.rom_rdata <= 32'h93804000;
          16'h1124 : blkif.rom_rdata <= 32'h1301c028;
          16'h1125 : blkif.rom_rdata <= 32'h23a02000;
          16'h1126 : blkif.rom_rdata <= 32'h9300f000;
          16'h1127 : blkif.rom_rdata <= 32'h33511000;
          16'h1128 : blkif.rom_rdata <= 32'h930e0000;
          16'h1129 : blkif.rom_rdata <= 32'h130ec028;
          16'h112a : blkif.rom_rdata <= 32'h6304d101;
          16'h112b : blkif.rom_rdata <= 32'h6f10002c;
          16'h112c : blkif.rom_rdata <= 32'hb7000080;
          16'h112d : blkif.rom_rdata <= 32'h93804000;
          16'h112e : blkif.rom_rdata <= 32'h1301d028;
          16'h112f : blkif.rom_rdata <= 32'h23a02000;
          16'h1130 : blkif.rom_rdata <= 32'h93000002;
          16'h1131 : blkif.rom_rdata <= 32'h33d10000;
          16'h1132 : blkif.rom_rdata <= 32'h930e0002;
          16'h1133 : blkif.rom_rdata <= 32'h130ed028;
          16'h1134 : blkif.rom_rdata <= 32'h6304d101;
          16'h1135 : blkif.rom_rdata <= 32'h6f108029;
          16'h1136 : blkif.rom_rdata <= 32'hb7000080;
          16'h1137 : blkif.rom_rdata <= 32'h93804000;
          16'h1138 : blkif.rom_rdata <= 32'h1301e028;
          16'h1139 : blkif.rom_rdata <= 32'h23a02000;
          16'h113a : blkif.rom_rdata <= 32'hb3500000;
          16'h113b : blkif.rom_rdata <= 32'h930e0000;
          16'h113c : blkif.rom_rdata <= 32'h130ee028;
          16'h113d : blkif.rom_rdata <= 32'h6384d001;
          16'h113e : blkif.rom_rdata <= 32'h6f104027;
          16'h113f : blkif.rom_rdata <= 32'hb7000080;
          16'h1140 : blkif.rom_rdata <= 32'h93804000;
          16'h1141 : blkif.rom_rdata <= 32'h1301f028;
          16'h1142 : blkif.rom_rdata <= 32'h23a02000;
          16'h1143 : blkif.rom_rdata <= 32'h93000040;
          16'h1144 : blkif.rom_rdata <= 32'h37110000;
          16'h1145 : blkif.rom_rdata <= 32'h13010180;
          16'h1146 : blkif.rom_rdata <= 32'h33d02000;
          16'h1147 : blkif.rom_rdata <= 32'h930e0000;
          16'h1148 : blkif.rom_rdata <= 32'h130ef028;
          16'h1149 : blkif.rom_rdata <= 32'h6304d001;
          16'h114a : blkif.rom_rdata <= 32'h6f104024;
          16'h114b : blkif.rom_rdata <= 32'hb7000080;
          16'h114c : blkif.rom_rdata <= 32'h93804000;
          16'h114d : blkif.rom_rdata <= 32'h13010029;
          16'h114e : blkif.rom_rdata <= 32'h23a02000;
          16'h114f : blkif.rom_rdata <= 32'hb780ffff;
          16'h1150 : blkif.rom_rdata <= 32'h93d10000;
          16'h1151 : blkif.rom_rdata <= 32'hb78effff;
          16'h1152 : blkif.rom_rdata <= 32'h130e0029;
          16'h1153 : blkif.rom_rdata <= 32'h6384d101;
          16'h1154 : blkif.rom_rdata <= 32'h6f10c021;
          16'h1155 : blkif.rom_rdata <= 32'hb7000080;
          16'h1156 : blkif.rom_rdata <= 32'h93804000;
          16'h1157 : blkif.rom_rdata <= 32'h13011029;
          16'h1158 : blkif.rom_rdata <= 32'h23a02000;
          16'h1159 : blkif.rom_rdata <= 32'hb780ffff;
          16'h115a : blkif.rom_rdata <= 32'h93d11000;
          16'h115b : blkif.rom_rdata <= 32'hb7ceff7f;
          16'h115c : blkif.rom_rdata <= 32'h130e1029;
          16'h115d : blkif.rom_rdata <= 32'h6384d101;
          16'h115e : blkif.rom_rdata <= 32'h6f10401f;
          16'h115f : blkif.rom_rdata <= 32'hb7000080;
          16'h1160 : blkif.rom_rdata <= 32'h93804000;
          16'h1161 : blkif.rom_rdata <= 32'h13015029;
          16'h1162 : blkif.rom_rdata <= 32'h23a02000;
          16'h1163 : blkif.rom_rdata <= 32'h9300f0ff;
          16'h1164 : blkif.rom_rdata <= 32'h93d10000;
          16'h1165 : blkif.rom_rdata <= 32'h930ef0ff;
          16'h1166 : blkif.rom_rdata <= 32'h130e5029;
          16'h1167 : blkif.rom_rdata <= 32'h6384d101;
          16'h1168 : blkif.rom_rdata <= 32'h6f10c01c;
          16'h1169 : blkif.rom_rdata <= 32'hb7000080;
          16'h116a : blkif.rom_rdata <= 32'h93804000;
          16'h116b : blkif.rom_rdata <= 32'h1301a029;
          16'h116c : blkif.rom_rdata <= 32'h23a02000;
          16'h116d : blkif.rom_rdata <= 32'hb7202121;
          16'h116e : blkif.rom_rdata <= 32'h93801012;
          16'h116f : blkif.rom_rdata <= 32'h93d10000;
          16'h1170 : blkif.rom_rdata <= 32'hb72e2121;
          16'h1171 : blkif.rom_rdata <= 32'h938e1e12;
          16'h1172 : blkif.rom_rdata <= 32'h130ea029;
          16'h1173 : blkif.rom_rdata <= 32'h6384d101;
          16'h1174 : blkif.rom_rdata <= 32'h6f10c019;
          16'h1175 : blkif.rom_rdata <= 32'hb7000080;
          16'h1176 : blkif.rom_rdata <= 32'h93804000;
          16'h1177 : blkif.rom_rdata <= 32'h1301f029;
          16'h1178 : blkif.rom_rdata <= 32'h23a02000;
          16'h1179 : blkif.rom_rdata <= 32'hb780ffff;
          16'h117a : blkif.rom_rdata <= 32'h93d01000;
          16'h117b : blkif.rom_rdata <= 32'hb7ceff7f;
          16'h117c : blkif.rom_rdata <= 32'h130ef029;
          16'h117d : blkif.rom_rdata <= 32'h6384d001;
          16'h117e : blkif.rom_rdata <= 32'h6f104017;
          16'h117f : blkif.rom_rdata <= 32'hb7000080;
          16'h1180 : blkif.rom_rdata <= 32'h93804000;
          16'h1181 : blkif.rom_rdata <= 32'h1301002a;
          16'h1182 : blkif.rom_rdata <= 32'h23a02000;
          16'h1183 : blkif.rom_rdata <= 32'h13020000;
          16'h1184 : blkif.rom_rdata <= 32'hb780ffff;
          16'h1185 : blkif.rom_rdata <= 32'h93d11000;
          16'h1186 : blkif.rom_rdata <= 32'h13830100;
          16'h1187 : blkif.rom_rdata <= 32'h13021200;
          16'h1188 : blkif.rom_rdata <= 32'h93022000;
          16'h1189 : blkif.rom_rdata <= 32'he31652fe;
          16'h118a : blkif.rom_rdata <= 32'hb7ceff7f;
          16'h118b : blkif.rom_rdata <= 32'h130e002a;
          16'h118c : blkif.rom_rdata <= 32'h6304d301;
          16'h118d : blkif.rom_rdata <= 32'h6f108013;
          16'h118e : blkif.rom_rdata <= 32'hb7000080;
          16'h118f : blkif.rom_rdata <= 32'h93804000;
          16'h1190 : blkif.rom_rdata <= 32'h1301302a;
          16'h1191 : blkif.rom_rdata <= 32'h23a02000;
          16'h1192 : blkif.rom_rdata <= 32'h13020000;
          16'h1193 : blkif.rom_rdata <= 32'hb780ffff;
          16'h1194 : blkif.rom_rdata <= 32'h93d11000;
          16'h1195 : blkif.rom_rdata <= 32'h13021200;
          16'h1196 : blkif.rom_rdata <= 32'h93022000;
          16'h1197 : blkif.rom_rdata <= 32'he31852fe;
          16'h1198 : blkif.rom_rdata <= 32'hb7ceff7f;
          16'h1199 : blkif.rom_rdata <= 32'h130e302a;
          16'h119a : blkif.rom_rdata <= 32'h6384d101;
          16'h119b : blkif.rom_rdata <= 32'h6f100010;
          16'h119c : blkif.rom_rdata <= 32'hb7000080;
          16'h119d : blkif.rom_rdata <= 32'h93804000;
          16'h119e : blkif.rom_rdata <= 32'h1301502a;
          16'h119f : blkif.rom_rdata <= 32'h23a02000;
          16'h11a0 : blkif.rom_rdata <= 32'h13020000;
          16'h11a1 : blkif.rom_rdata <= 32'hb780ffff;
          16'h11a2 : blkif.rom_rdata <= 32'h13000000;
          16'h11a3 : blkif.rom_rdata <= 32'h13000000;
          16'h11a4 : blkif.rom_rdata <= 32'h93d1f000;
          16'h11a5 : blkif.rom_rdata <= 32'h13021200;
          16'h11a6 : blkif.rom_rdata <= 32'h93022000;
          16'h11a7 : blkif.rom_rdata <= 32'he31452fe;
          16'h11a8 : blkif.rom_rdata <= 32'hb70e0200;
          16'h11a9 : blkif.rom_rdata <= 32'h938efeff;
          16'h11aa : blkif.rom_rdata <= 32'h130e502a;
          16'h11ab : blkif.rom_rdata <= 32'h6384d101;
          16'h11ac : blkif.rom_rdata <= 32'h6f10c00b;
          16'h11ad : blkif.rom_rdata <= 32'hb7000080;
          16'h11ae : blkif.rom_rdata <= 32'h93804000;
          16'h11af : blkif.rom_rdata <= 32'h1301602a;
          16'h11b0 : blkif.rom_rdata <= 32'h23a02000;
          16'h11b1 : blkif.rom_rdata <= 32'h9350f001;
          16'h11b2 : blkif.rom_rdata <= 32'h930e0000;
          16'h11b3 : blkif.rom_rdata <= 32'h130e602a;
          16'h11b4 : blkif.rom_rdata <= 32'h6384d001;
          16'h11b5 : blkif.rom_rdata <= 32'h6f108009;
          16'h11b6 : blkif.rom_rdata <= 32'hb7000080;
          16'h11b7 : blkif.rom_rdata <= 32'h93804000;
          16'h11b8 : blkif.rom_rdata <= 32'h1301702a;
          16'h11b9 : blkif.rom_rdata <= 32'h23a02000;
          16'h11ba : blkif.rom_rdata <= 32'h93001002;
          16'h11bb : blkif.rom_rdata <= 32'h13d04001;
          16'h11bc : blkif.rom_rdata <= 32'h930e0000;
          16'h11bd : blkif.rom_rdata <= 32'h130e702a;
          16'h11be : blkif.rom_rdata <= 32'h6304d001;
          16'h11bf : blkif.rom_rdata <= 32'h6f100007;
          16'h11c0 : blkif.rom_rdata <= 32'hb7000080;
          16'h11c1 : blkif.rom_rdata <= 32'h93804000;
          16'h11c2 : blkif.rom_rdata <= 32'h1301802a;
          16'h11c3 : blkif.rom_rdata <= 32'h23a02000;
          16'h11c4 : blkif.rom_rdata <= 32'h93000000;
          16'h11c5 : blkif.rom_rdata <= 32'h13010000;
          16'h11c6 : blkif.rom_rdata <= 32'hb3812040;
          16'h11c7 : blkif.rom_rdata <= 32'h930e0000;
          16'h11c8 : blkif.rom_rdata <= 32'h130e802a;
          16'h11c9 : blkif.rom_rdata <= 32'h6384d101;
          16'h11ca : blkif.rom_rdata <= 32'h6f104004;
          16'h11cb : blkif.rom_rdata <= 32'hb7000080;
          16'h11cc : blkif.rom_rdata <= 32'h93804000;
          16'h11cd : blkif.rom_rdata <= 32'h1301a02a;
          16'h11ce : blkif.rom_rdata <= 32'h23a02000;
          16'h11cf : blkif.rom_rdata <= 32'h93003000;
          16'h11d0 : blkif.rom_rdata <= 32'h13017000;
          16'h11d1 : blkif.rom_rdata <= 32'hb3812040;
          16'h11d2 : blkif.rom_rdata <= 32'h930ec0ff;
          16'h11d3 : blkif.rom_rdata <= 32'h130ea02a;
          16'h11d4 : blkif.rom_rdata <= 32'h6384d101;
          16'h11d5 : blkif.rom_rdata <= 32'h6f108001;
          16'h11d6 : blkif.rom_rdata <= 32'hb7000080;
          16'h11d7 : blkif.rom_rdata <= 32'h93804000;
          16'h11d8 : blkif.rom_rdata <= 32'h1301302b;
          16'h11d9 : blkif.rom_rdata <= 32'h23a02000;
          16'h11da : blkif.rom_rdata <= 32'h93000000;
          16'h11db : blkif.rom_rdata <= 32'h1301f0ff;
          16'h11dc : blkif.rom_rdata <= 32'hb3812040;
          16'h11dd : blkif.rom_rdata <= 32'h930e1000;
          16'h11de : blkif.rom_rdata <= 32'h130e302b;
          16'h11df : blkif.rom_rdata <= 32'he398d17f;
          16'h11e0 : blkif.rom_rdata <= 32'hb7000080;
          16'h11e1 : blkif.rom_rdata <= 32'h93804000;
          16'h11e2 : blkif.rom_rdata <= 32'h1301502b;
          16'h11e3 : blkif.rom_rdata <= 32'h23a02000;
          16'h11e4 : blkif.rom_rdata <= 32'h9300f0ff;
          16'h11e5 : blkif.rom_rdata <= 32'h1301f0ff;
          16'h11e6 : blkif.rom_rdata <= 32'hb3812040;
          16'h11e7 : blkif.rom_rdata <= 32'h930e0000;
          16'h11e8 : blkif.rom_rdata <= 32'h130e502b;
          16'h11e9 : blkif.rom_rdata <= 32'he394d17d;
          16'h11ea : blkif.rom_rdata <= 32'hb7000080;
          16'h11eb : blkif.rom_rdata <= 32'h93804000;
          16'h11ec : blkif.rom_rdata <= 32'h1301602b;
          16'h11ed : blkif.rom_rdata <= 32'h23a02000;
          16'h11ee : blkif.rom_rdata <= 32'h9300d000;
          16'h11ef : blkif.rom_rdata <= 32'h1301b000;
          16'h11f0 : blkif.rom_rdata <= 32'hb3802040;
          16'h11f1 : blkif.rom_rdata <= 32'h930e2000;
          16'h11f2 : blkif.rom_rdata <= 32'h130e602b;
          16'h11f3 : blkif.rom_rdata <= 32'he390d07b;
          16'h11f4 : blkif.rom_rdata <= 32'hb7000080;
          16'h11f5 : blkif.rom_rdata <= 32'h93804000;
          16'h11f6 : blkif.rom_rdata <= 32'h1301702b;
          16'h11f7 : blkif.rom_rdata <= 32'h23a02000;
          16'h11f8 : blkif.rom_rdata <= 32'h9300e000;
          16'h11f9 : blkif.rom_rdata <= 32'h1301b000;
          16'h11fa : blkif.rom_rdata <= 32'h33812040;
          16'h11fb : blkif.rom_rdata <= 32'h930e3000;
          16'h11fc : blkif.rom_rdata <= 32'h130e702b;
          16'h11fd : blkif.rom_rdata <= 32'he31cd177;
          16'h11fe : blkif.rom_rdata <= 32'hb7000080;
          16'h11ff : blkif.rom_rdata <= 32'h93804000;
          16'h1200 : blkif.rom_rdata <= 32'h1301802b;
          16'h1201 : blkif.rom_rdata <= 32'h23a02000;
          16'h1202 : blkif.rom_rdata <= 32'h9300d000;
          16'h1203 : blkif.rom_rdata <= 32'hb3801040;
          16'h1204 : blkif.rom_rdata <= 32'h930e0000;
          16'h1205 : blkif.rom_rdata <= 32'h130e802b;
          16'h1206 : blkif.rom_rdata <= 32'he39ad075;
          16'h1207 : blkif.rom_rdata <= 32'hb7000080;
          16'h1208 : blkif.rom_rdata <= 32'h93804000;
          16'h1209 : blkif.rom_rdata <= 32'h1301902b;
          16'h120a : blkif.rom_rdata <= 32'h23a02000;
          16'h120b : blkif.rom_rdata <= 32'h13020000;
          16'h120c : blkif.rom_rdata <= 32'h9300d000;
          16'h120d : blkif.rom_rdata <= 32'h1301b000;
          16'h120e : blkif.rom_rdata <= 32'hb3812040;
          16'h120f : blkif.rom_rdata <= 32'h13830100;
          16'h1210 : blkif.rom_rdata <= 32'h13021200;
          16'h1211 : blkif.rom_rdata <= 32'h93022000;
          16'h1212 : blkif.rom_rdata <= 32'he31452fe;
          16'h1213 : blkif.rom_rdata <= 32'h930e2000;
          16'h1214 : blkif.rom_rdata <= 32'h130e902b;
          16'h1215 : blkif.rom_rdata <= 32'he31cd371;
          16'h1216 : blkif.rom_rdata <= 32'hb7000080;
          16'h1217 : blkif.rom_rdata <= 32'h93804000;
          16'h1218 : blkif.rom_rdata <= 32'h1301c02b;
          16'h1219 : blkif.rom_rdata <= 32'h23a02000;
          16'h121a : blkif.rom_rdata <= 32'h13020000;
          16'h121b : blkif.rom_rdata <= 32'h9300d000;
          16'h121c : blkif.rom_rdata <= 32'h1301b000;
          16'h121d : blkif.rom_rdata <= 32'hb3812040;
          16'h121e : blkif.rom_rdata <= 32'h13021200;
          16'h121f : blkif.rom_rdata <= 32'h93022000;
          16'h1220 : blkif.rom_rdata <= 32'he31652fe;
          16'h1221 : blkif.rom_rdata <= 32'h930e2000;
          16'h1222 : blkif.rom_rdata <= 32'h130ec02b;
          16'h1223 : blkif.rom_rdata <= 32'he390d16f;
          16'h1224 : blkif.rom_rdata <= 32'hb7000080;
          16'h1225 : blkif.rom_rdata <= 32'h93804000;
          16'h1226 : blkif.rom_rdata <= 32'h1301102c;
          16'h1227 : blkif.rom_rdata <= 32'h23a02000;
          16'h1228 : blkif.rom_rdata <= 32'h13020000;
          16'h1229 : blkif.rom_rdata <= 32'h9300f000;
          16'h122a : blkif.rom_rdata <= 32'h13000000;
          16'h122b : blkif.rom_rdata <= 32'h13000000;
          16'h122c : blkif.rom_rdata <= 32'h1301b000;
          16'h122d : blkif.rom_rdata <= 32'hb3812040;
          16'h122e : blkif.rom_rdata <= 32'h13021200;
          16'h122f : blkif.rom_rdata <= 32'h93022000;
          16'h1230 : blkif.rom_rdata <= 32'he31252fe;
          16'h1231 : blkif.rom_rdata <= 32'h930e4000;
          16'h1232 : blkif.rom_rdata <= 32'h130e102c;
          16'h1233 : blkif.rom_rdata <= 32'he390d16b;
          16'h1234 : blkif.rom_rdata <= 32'hb7000080;
          16'h1235 : blkif.rom_rdata <= 32'h93804000;
          16'h1236 : blkif.rom_rdata <= 32'h1301202c;
          16'h1237 : blkif.rom_rdata <= 32'h23a02000;
          16'h1238 : blkif.rom_rdata <= 32'h13020000;
          16'h1239 : blkif.rom_rdata <= 32'h1301b000;
          16'h123a : blkif.rom_rdata <= 32'h9300d000;
          16'h123b : blkif.rom_rdata <= 32'hb3812040;
          16'h123c : blkif.rom_rdata <= 32'h13021200;
          16'h123d : blkif.rom_rdata <= 32'h93022000;
          16'h123e : blkif.rom_rdata <= 32'he31652fe;
          16'h123f : blkif.rom_rdata <= 32'h930e2000;
          16'h1240 : blkif.rom_rdata <= 32'h130e202c;
          16'h1241 : blkif.rom_rdata <= 32'he394d167;
          16'h1242 : blkif.rom_rdata <= 32'hb7000080;
          16'h1243 : blkif.rom_rdata <= 32'h93804000;
          16'h1244 : blkif.rom_rdata <= 32'h1301402c;
          16'h1245 : blkif.rom_rdata <= 32'h23a02000;
          16'h1246 : blkif.rom_rdata <= 32'h13020000;
          16'h1247 : blkif.rom_rdata <= 32'h1301b000;
          16'h1248 : blkif.rom_rdata <= 32'h9300f000;
          16'h1249 : blkif.rom_rdata <= 32'h13000000;
          16'h124a : blkif.rom_rdata <= 32'h13000000;
          16'h124b : blkif.rom_rdata <= 32'hb3812040;
          16'h124c : blkif.rom_rdata <= 32'h13021200;
          16'h124d : blkif.rom_rdata <= 32'h93022000;
          16'h124e : blkif.rom_rdata <= 32'he31252fe;
          16'h124f : blkif.rom_rdata <= 32'h930e4000;
          16'h1250 : blkif.rom_rdata <= 32'h130e402c;
          16'h1251 : blkif.rom_rdata <= 32'he394d163;
          16'h1252 : blkif.rom_rdata <= 32'hb7000080;
          16'h1253 : blkif.rom_rdata <= 32'h93804000;
          16'h1254 : blkif.rom_rdata <= 32'h1301802c;
          16'h1255 : blkif.rom_rdata <= 32'h23a02000;
          16'h1256 : blkif.rom_rdata <= 32'h930010ff;
          16'h1257 : blkif.rom_rdata <= 32'h33011040;
          16'h1258 : blkif.rom_rdata <= 32'h930ef000;
          16'h1259 : blkif.rom_rdata <= 32'h130e802c;
          16'h125a : blkif.rom_rdata <= 32'he312d161;
          16'h125b : blkif.rom_rdata <= 32'hb7000080;
          16'h125c : blkif.rom_rdata <= 32'h93804000;
          16'h125d : blkif.rom_rdata <= 32'h1301902c;
          16'h125e : blkif.rom_rdata <= 32'h23a02000;
          16'h125f : blkif.rom_rdata <= 32'h93000002;
          16'h1260 : blkif.rom_rdata <= 32'h33810040;
          16'h1261 : blkif.rom_rdata <= 32'h930e0002;
          16'h1262 : blkif.rom_rdata <= 32'h130e902c;
          16'h1263 : blkif.rom_rdata <= 32'he310d15f;
          16'h1264 : blkif.rom_rdata <= 32'hb7000080;
          16'h1265 : blkif.rom_rdata <= 32'h93804000;
          16'h1266 : blkif.rom_rdata <= 32'h1301a02c;
          16'h1267 : blkif.rom_rdata <= 32'h23a02000;
          16'h1268 : blkif.rom_rdata <= 32'hb3000040;
          16'h1269 : blkif.rom_rdata <= 32'h930e0000;
          16'h126a : blkif.rom_rdata <= 32'h130ea02c;
          16'h126b : blkif.rom_rdata <= 32'he390d05d;
          16'h126c : blkif.rom_rdata <= 32'hb7000080;
          16'h126d : blkif.rom_rdata <= 32'h93804000;
          16'h126e : blkif.rom_rdata <= 32'h1301b02c;
          16'h126f : blkif.rom_rdata <= 32'h23a02000;
          16'h1270 : blkif.rom_rdata <= 32'h93000001;
          16'h1271 : blkif.rom_rdata <= 32'h1301e001;
          16'h1272 : blkif.rom_rdata <= 32'h33802040;
          16'h1273 : blkif.rom_rdata <= 32'h930e0000;
          16'h1274 : blkif.rom_rdata <= 32'h130eb02c;
          16'h1275 : blkif.rom_rdata <= 32'he31cd059;
          16'h1276 : blkif.rom_rdata <= 32'hb7000080;
          16'h1277 : blkif.rom_rdata <= 32'h93804000;
          16'h1278 : blkif.rom_rdata <= 32'h1301c02c;
          16'h1279 : blkif.rom_rdata <= 32'h23a02000;
          16'h127a : blkif.rom_rdata <= 32'h97300000;
          16'h127b : blkif.rom_rdata <= 32'h93808064;
          16'h127c : blkif.rom_rdata <= 32'h3701aa00;
          16'h127d : blkif.rom_rdata <= 32'h1301a10a;
          16'h127e : blkif.rom_rdata <= 32'h23a02000;
          16'h127f : blkif.rom_rdata <= 32'h83a10000;
          16'h1280 : blkif.rom_rdata <= 32'hb70eaa00;
          16'h1281 : blkif.rom_rdata <= 32'h938eae0a;
          16'h1282 : blkif.rom_rdata <= 32'h130ec02c;
          16'h1283 : blkif.rom_rdata <= 32'he390d157;
          16'h1284 : blkif.rom_rdata <= 32'hb7000080;
          16'h1285 : blkif.rom_rdata <= 32'h93804000;
          16'h1286 : blkif.rom_rdata <= 32'h1301f02c;
          16'h1287 : blkif.rom_rdata <= 32'h23a02000;
          16'h1288 : blkif.rom_rdata <= 32'h97300000;
          16'h1289 : blkif.rom_rdata <= 32'h93800061;
          16'h128a : blkif.rom_rdata <= 32'h37a10aa0;
          16'h128b : blkif.rom_rdata <= 32'h1301a100;
          16'h128c : blkif.rom_rdata <= 32'h23a62000;
          16'h128d : blkif.rom_rdata <= 32'h83a1c000;
          16'h128e : blkif.rom_rdata <= 32'hb7ae0aa0;
          16'h128f : blkif.rom_rdata <= 32'h938eae00;
          16'h1290 : blkif.rom_rdata <= 32'h130ef02c;
          16'h1291 : blkif.rom_rdata <= 32'he394d153;
          16'h1292 : blkif.rom_rdata <= 32'hb7000080;
          16'h1293 : blkif.rom_rdata <= 32'h93804000;
          16'h1294 : blkif.rom_rdata <= 32'h1301002d;
          16'h1295 : blkif.rom_rdata <= 32'h23a02000;
          16'h1296 : blkif.rom_rdata <= 32'h97300000;
          16'h1297 : blkif.rom_rdata <= 32'h9380405f;
          16'h1298 : blkif.rom_rdata <= 32'h3701aa00;
          16'h1299 : blkif.rom_rdata <= 32'h1301a10a;
          16'h129a : blkif.rom_rdata <= 32'h23aa20fe;
          16'h129b : blkif.rom_rdata <= 32'h83a140ff;
          16'h129c : blkif.rom_rdata <= 32'hb70eaa00;
          16'h129d : blkif.rom_rdata <= 32'h938eae0a;
          16'h129e : blkif.rom_rdata <= 32'h130e002d;
          16'h129f : blkif.rom_rdata <= 32'he398d14f;
          16'h12a0 : blkif.rom_rdata <= 32'hb7000080;
          16'h12a1 : blkif.rom_rdata <= 32'h93804000;
          16'h12a2 : blkif.rom_rdata <= 32'h1301102d;
          16'h12a3 : blkif.rom_rdata <= 32'h23a02000;
          16'h12a4 : blkif.rom_rdata <= 32'h97300000;
          16'h12a5 : blkif.rom_rdata <= 32'h9380c05b;
          16'h12a6 : blkif.rom_rdata <= 32'h37b100aa;
          16'h12a7 : blkif.rom_rdata <= 32'h130101a0;
          16'h12a8 : blkif.rom_rdata <= 32'h23ac20fe;
          16'h12a9 : blkif.rom_rdata <= 32'h83a180ff;
          16'h12aa : blkif.rom_rdata <= 32'hb7be00aa;
          16'h12ab : blkif.rom_rdata <= 32'h938e0ea0;
          16'h12ac : blkif.rom_rdata <= 32'h130e102d;
          16'h12ad : blkif.rom_rdata <= 32'he39cd14b;
          16'h12ae : blkif.rom_rdata <= 32'hb7000080;
          16'h12af : blkif.rom_rdata <= 32'h93804000;
          16'h12b0 : blkif.rom_rdata <= 32'h1301402d;
          16'h12b1 : blkif.rom_rdata <= 32'h23a02000;
          16'h12b2 : blkif.rom_rdata <= 32'h97300000;
          16'h12b3 : blkif.rom_rdata <= 32'h93808058;
          16'h12b4 : blkif.rom_rdata <= 32'h37513412;
          16'h12b5 : blkif.rom_rdata <= 32'h13018167;
          16'h12b6 : blkif.rom_rdata <= 32'h138200fe;
          16'h12b7 : blkif.rom_rdata <= 32'h23202202;
          16'h12b8 : blkif.rom_rdata <= 32'h83a10000;
          16'h12b9 : blkif.rom_rdata <= 32'hb75e3412;
          16'h12ba : blkif.rom_rdata <= 32'h938e8e67;
          16'h12bb : blkif.rom_rdata <= 32'h130e402d;
          16'h12bc : blkif.rom_rdata <= 32'he39ed147;
          16'h12bd : blkif.rom_rdata <= 32'hb7000080;
          16'h12be : blkif.rom_rdata <= 32'h93804000;
          16'h12bf : blkif.rom_rdata <= 32'h1301502d;
          16'h12c0 : blkif.rom_rdata <= 32'h23a02000;
          16'h12c1 : blkif.rom_rdata <= 32'h97300000;
          16'h12c2 : blkif.rom_rdata <= 32'h9380c054;
          16'h12c3 : blkif.rom_rdata <= 32'h37312158;
          16'h12c4 : blkif.rom_rdata <= 32'h13018109;
          16'h12c5 : blkif.rom_rdata <= 32'h9380d0ff;
          16'h12c6 : blkif.rom_rdata <= 32'ha3a32000;
          16'h12c7 : blkif.rom_rdata <= 32'h17320000;
          16'h12c8 : blkif.rom_rdata <= 32'h13028253;
          16'h12c9 : blkif.rom_rdata <= 32'h83210200;
          16'h12ca : blkif.rom_rdata <= 32'hb73e2158;
          16'h12cb : blkif.rom_rdata <= 32'h938e8e09;
          16'h12cc : blkif.rom_rdata <= 32'h130e502d;
          16'h12cd : blkif.rom_rdata <= 32'he39cd143;
          16'h12ce : blkif.rom_rdata <= 32'h130e602d;
          16'h12cf : blkif.rom_rdata <= 32'h13020000;
          16'h12d0 : blkif.rom_rdata <= 32'hb7d0bbaa;
          16'h12d1 : blkif.rom_rdata <= 32'h9380d0cd;
          16'h12d2 : blkif.rom_rdata <= 32'h17310000;
          16'h12d3 : blkif.rom_rdata <= 32'h1301814e;
          16'h12d4 : blkif.rom_rdata <= 32'h23201100;
          16'h12d5 : blkif.rom_rdata <= 32'h83210100;
          16'h12d6 : blkif.rom_rdata <= 32'hb7debbaa;
          16'h12d7 : blkif.rom_rdata <= 32'h938edecd;
          16'h12d8 : blkif.rom_rdata <= 32'he396d141;
          16'h12d9 : blkif.rom_rdata <= 32'h13021200;
          16'h12da : blkif.rom_rdata <= 32'h93022000;
          16'h12db : blkif.rom_rdata <= 32'he31a52fc;
          16'h12dc : blkif.rom_rdata <= 32'h130eb02d;
          16'h12dd : blkif.rom_rdata <= 32'h13020000;
          16'h12de : blkif.rom_rdata <= 32'hb7e0cdbc;
          16'h12df : blkif.rom_rdata <= 32'h9380b0aa;
          16'h12e0 : blkif.rom_rdata <= 32'h13000000;
          16'h12e1 : blkif.rom_rdata <= 32'h13000000;
          16'h12e2 : blkif.rom_rdata <= 32'h17310000;
          16'h12e3 : blkif.rom_rdata <= 32'h1301814a;
          16'h12e4 : blkif.rom_rdata <= 32'h232a1100;
          16'h12e5 : blkif.rom_rdata <= 32'h83214101;
          16'h12e6 : blkif.rom_rdata <= 32'hb7eecdbc;
          16'h12e7 : blkif.rom_rdata <= 32'h938ebeaa;
          16'h12e8 : blkif.rom_rdata <= 32'he396d13d;
          16'h12e9 : blkif.rom_rdata <= 32'h13021200;
          16'h12ea : blkif.rom_rdata <= 32'h93022000;
          16'h12eb : blkif.rom_rdata <= 32'he31652fc;
          16'h12ec : blkif.rom_rdata <= 32'h130ec02d;
          16'h12ed : blkif.rom_rdata <= 32'h13020000;
          16'h12ee : blkif.rom_rdata <= 32'h17310000;
          16'h12ef : blkif.rom_rdata <= 32'h13018147;
          16'h12f0 : blkif.rom_rdata <= 32'hb7201100;
          16'h12f1 : blkif.rom_rdata <= 32'h93803023;
          16'h12f2 : blkif.rom_rdata <= 32'h23201100;
          16'h12f3 : blkif.rom_rdata <= 32'h83210100;
          16'h12f4 : blkif.rom_rdata <= 32'hb72e1100;
          16'h12f5 : blkif.rom_rdata <= 32'h938e3e23;
          16'h12f6 : blkif.rom_rdata <= 32'he39ad139;
          16'h12f7 : blkif.rom_rdata <= 32'h13021200;
          16'h12f8 : blkif.rom_rdata <= 32'h93022000;
          16'h12f9 : blkif.rom_rdata <= 32'he31a52fc;
          16'h12fa : blkif.rom_rdata <= 32'h130e102e;
          16'h12fb : blkif.rom_rdata <= 32'h13020000;
          16'h12fc : blkif.rom_rdata <= 32'h17310000;
          16'h12fd : blkif.rom_rdata <= 32'h13010144;
          16'h12fe : blkif.rom_rdata <= 32'h13000000;
          16'h12ff : blkif.rom_rdata <= 32'h13000000;
          16'h1300 : blkif.rom_rdata <= 32'hb7302312;
          16'h1301 : blkif.rom_rdata <= 32'h93801000;
          16'h1302 : blkif.rom_rdata <= 32'h232a1100;
          16'h1303 : blkif.rom_rdata <= 32'h83214101;
          16'h1304 : blkif.rom_rdata <= 32'hb73e2312;
          16'h1305 : blkif.rom_rdata <= 32'h938e1e00;
          16'h1306 : blkif.rom_rdata <= 32'he39ad135;
          16'h1307 : blkif.rom_rdata <= 32'h13021200;
          16'h1308 : blkif.rom_rdata <= 32'h93022000;
          16'h1309 : blkif.rom_rdata <= 32'he31652fc;
          16'h130a : blkif.rom_rdata <= 32'hb7000080;
          16'h130b : blkif.rom_rdata <= 32'h93804000;
          16'h130c : blkif.rom_rdata <= 32'h1301202e;
          16'h130d : blkif.rom_rdata <= 32'h23a02000;
          16'h130e : blkif.rom_rdata <= 32'hb70001ff;
          16'h130f : blkif.rom_rdata <= 32'h938000f0;
          16'h1310 : blkif.rom_rdata <= 32'h37110f0f;
          16'h1311 : blkif.rom_rdata <= 32'h1301f1f0;
          16'h1312 : blkif.rom_rdata <= 32'hb3c12000;
          16'h1313 : blkif.rom_rdata <= 32'hb7fe0ff0;
          16'h1314 : blkif.rom_rdata <= 32'h938efe00;
          16'h1315 : blkif.rom_rdata <= 32'h130e202e;
          16'h1316 : blkif.rom_rdata <= 32'he39ad131;
          16'h1317 : blkif.rom_rdata <= 32'hb7000080;
          16'h1318 : blkif.rom_rdata <= 32'h93804000;
          16'h1319 : blkif.rom_rdata <= 32'h1301502e;
          16'h131a : blkif.rom_rdata <= 32'h23a02000;
          16'h131b : blkif.rom_rdata <= 32'hb7f00ff0;
          16'h131c : blkif.rom_rdata <= 32'h9380f000;
          16'h131d : blkif.rom_rdata <= 32'h37f1f0f0;
          16'h131e : blkif.rom_rdata <= 32'h1301010f;
          16'h131f : blkif.rom_rdata <= 32'hb3c12000;
          16'h1320 : blkif.rom_rdata <= 32'hb70eff00;
          16'h1321 : blkif.rom_rdata <= 32'h938efe0f;
          16'h1322 : blkif.rom_rdata <= 32'h130e502e;
          16'h1323 : blkif.rom_rdata <= 32'he390d12f;
          16'h1324 : blkif.rom_rdata <= 32'hb7000080;
          16'h1325 : blkif.rom_rdata <= 32'h93804000;
          16'h1326 : blkif.rom_rdata <= 32'h1301602e;
          16'h1327 : blkif.rom_rdata <= 32'h23a02000;
          16'h1328 : blkif.rom_rdata <= 32'hb70001ff;
          16'h1329 : blkif.rom_rdata <= 32'h938000f0;
          16'h132a : blkif.rom_rdata <= 32'h37110f0f;
          16'h132b : blkif.rom_rdata <= 32'h1301f1f0;
          16'h132c : blkif.rom_rdata <= 32'hb3c02000;
          16'h132d : blkif.rom_rdata <= 32'hb7fe0ff0;
          16'h132e : blkif.rom_rdata <= 32'h938efe00;
          16'h132f : blkif.rom_rdata <= 32'h130e602e;
          16'h1330 : blkif.rom_rdata <= 32'he396d02b;
          16'h1331 : blkif.rom_rdata <= 32'hb7000080;
          16'h1332 : blkif.rom_rdata <= 32'h93804000;
          16'h1333 : blkif.rom_rdata <= 32'h1301702e;
          16'h1334 : blkif.rom_rdata <= 32'h23a02000;
          16'h1335 : blkif.rom_rdata <= 32'hb70001ff;
          16'h1336 : blkif.rom_rdata <= 32'h938000f0;
          16'h1337 : blkif.rom_rdata <= 32'h37110f0f;
          16'h1338 : blkif.rom_rdata <= 32'h1301f1f0;
          16'h1339 : blkif.rom_rdata <= 32'h33c12000;
          16'h133a : blkif.rom_rdata <= 32'hb7fe0ff0;
          16'h133b : blkif.rom_rdata <= 32'h938efe00;
          16'h133c : blkif.rom_rdata <= 32'h130e702e;
          16'h133d : blkif.rom_rdata <= 32'he31cd127;
          16'h133e : blkif.rom_rdata <= 32'hb7000080;
          16'h133f : blkif.rom_rdata <= 32'h93804000;
          16'h1340 : blkif.rom_rdata <= 32'h1301802e;
          16'h1341 : blkif.rom_rdata <= 32'h23a02000;
          16'h1342 : blkif.rom_rdata <= 32'hb70001ff;
          16'h1343 : blkif.rom_rdata <= 32'h938000f0;
          16'h1344 : blkif.rom_rdata <= 32'hb3c01000;
          16'h1345 : blkif.rom_rdata <= 32'h930e0000;
          16'h1346 : blkif.rom_rdata <= 32'h130e802e;
          16'h1347 : blkif.rom_rdata <= 32'he398d025;
          16'h1348 : blkif.rom_rdata <= 32'hb7000080;
          16'h1349 : blkif.rom_rdata <= 32'h93804000;
          16'h134a : blkif.rom_rdata <= 32'h1301902e;
          16'h134b : blkif.rom_rdata <= 32'h23a02000;
          16'h134c : blkif.rom_rdata <= 32'h13020000;
          16'h134d : blkif.rom_rdata <= 32'hb70001ff;
          16'h134e : blkif.rom_rdata <= 32'h938000f0;
          16'h134f : blkif.rom_rdata <= 32'h37110f0f;
          16'h1350 : blkif.rom_rdata <= 32'h1301f1f0;
          16'h1351 : blkif.rom_rdata <= 32'hb3c12000;
          16'h1352 : blkif.rom_rdata <= 32'h13830100;
          16'h1353 : blkif.rom_rdata <= 32'h13021200;
          16'h1354 : blkif.rom_rdata <= 32'h93022000;
          16'h1355 : blkif.rom_rdata <= 32'he31052fe;
          16'h1356 : blkif.rom_rdata <= 32'hb7fe0ff0;
          16'h1357 : blkif.rom_rdata <= 32'h938efe00;
          16'h1358 : blkif.rom_rdata <= 32'h130e902e;
          16'h1359 : blkif.rom_rdata <= 32'he314d321;
          16'h135a : blkif.rom_rdata <= 32'hb7000080;
          16'h135b : blkif.rom_rdata <= 32'h93804000;
          16'h135c : blkif.rom_rdata <= 32'h1301a02e;
          16'h135d : blkif.rom_rdata <= 32'h23a02000;
          16'h135e : blkif.rom_rdata <= 32'h13020000;
          16'h135f : blkif.rom_rdata <= 32'hb710f00f;
          16'h1360 : blkif.rom_rdata <= 32'h938000ff;
          16'h1361 : blkif.rom_rdata <= 32'h37f1f0f0;
          16'h1362 : blkif.rom_rdata <= 32'h1301010f;
          16'h1363 : blkif.rom_rdata <= 32'hb3c12000;
          16'h1364 : blkif.rom_rdata <= 32'h13000000;
          16'h1365 : blkif.rom_rdata <= 32'h13830100;
          16'h1366 : blkif.rom_rdata <= 32'h13021200;
          16'h1367 : blkif.rom_rdata <= 32'h93022000;
          16'h1368 : blkif.rom_rdata <= 32'he31e52fc;
          16'h1369 : blkif.rom_rdata <= 32'hb70e01ff;
          16'h136a : blkif.rom_rdata <= 32'h938e0ef0;
          16'h136b : blkif.rom_rdata <= 32'h130ea02e;
          16'h136c : blkif.rom_rdata <= 32'he31ed31b;
          16'h136d : blkif.rom_rdata <= 32'hb7000080;
          16'h136e : blkif.rom_rdata <= 32'h93804000;
          16'h136f : blkif.rom_rdata <= 32'h1301c02e;
          16'h1370 : blkif.rom_rdata <= 32'h23a02000;
          16'h1371 : blkif.rom_rdata <= 32'h13020000;
          16'h1372 : blkif.rom_rdata <= 32'hb70001ff;
          16'h1373 : blkif.rom_rdata <= 32'h938000f0;
          16'h1374 : blkif.rom_rdata <= 32'h37110f0f;
          16'h1375 : blkif.rom_rdata <= 32'h1301f1f0;
          16'h1376 : blkif.rom_rdata <= 32'hb3c12000;
          16'h1377 : blkif.rom_rdata <= 32'h13021200;
          16'h1378 : blkif.rom_rdata <= 32'h93022000;
          16'h1379 : blkif.rom_rdata <= 32'he31252fe;
          16'h137a : blkif.rom_rdata <= 32'hb7fe0ff0;
          16'h137b : blkif.rom_rdata <= 32'h938efe00;
          16'h137c : blkif.rom_rdata <= 32'h130ec02e;
          16'h137d : blkif.rom_rdata <= 32'he39cd117;
          16'h137e : blkif.rom_rdata <= 32'hb7000080;
          16'h137f : blkif.rom_rdata <= 32'h93804000;
          16'h1380 : blkif.rom_rdata <= 32'h1301102f;
          16'h1381 : blkif.rom_rdata <= 32'h23a02000;
          16'h1382 : blkif.rom_rdata <= 32'h13020000;
          16'h1383 : blkif.rom_rdata <= 32'hb700ff00;
          16'h1384 : blkif.rom_rdata <= 32'h9380f00f;
          16'h1385 : blkif.rom_rdata <= 32'h13000000;
          16'h1386 : blkif.rom_rdata <= 32'h13000000;
          16'h1387 : blkif.rom_rdata <= 32'h37110f0f;
          16'h1388 : blkif.rom_rdata <= 32'h1301f1f0;
          16'h1389 : blkif.rom_rdata <= 32'hb3c12000;
          16'h138a : blkif.rom_rdata <= 32'h13021200;
          16'h138b : blkif.rom_rdata <= 32'h93022000;
          16'h138c : blkif.rom_rdata <= 32'he31e52fc;
          16'h138d : blkif.rom_rdata <= 32'hb71ef00f;
          16'h138e : blkif.rom_rdata <= 32'h938e0eff;
          16'h138f : blkif.rom_rdata <= 32'h130e102f;
          16'h1390 : blkif.rom_rdata <= 32'he396d113;
          16'h1391 : blkif.rom_rdata <= 32'hb7000080;
          16'h1392 : blkif.rom_rdata <= 32'h93804000;
          16'h1393 : blkif.rom_rdata <= 32'h1301802f;
          16'h1394 : blkif.rom_rdata <= 32'h23a02000;
          16'h1395 : blkif.rom_rdata <= 32'hb70001ff;
          16'h1396 : blkif.rom_rdata <= 32'h938000f0;
          16'h1397 : blkif.rom_rdata <= 32'h33411000;
          16'h1398 : blkif.rom_rdata <= 32'hb70e01ff;
          16'h1399 : blkif.rom_rdata <= 32'h938e0ef0;
          16'h139a : blkif.rom_rdata <= 32'h130e802f;
          16'h139b : blkif.rom_rdata <= 32'he310d111;
          16'h139c : blkif.rom_rdata <= 32'hb7000080;
          16'h139d : blkif.rom_rdata <= 32'h93804000;
          16'h139e : blkif.rom_rdata <= 32'h1301902f;
          16'h139f : blkif.rom_rdata <= 32'h23a02000;
          16'h13a0 : blkif.rom_rdata <= 32'hb700ff00;
          16'h13a1 : blkif.rom_rdata <= 32'h9380f00f;
          16'h13a2 : blkif.rom_rdata <= 32'h33c10000;
          16'h13a3 : blkif.rom_rdata <= 32'hb70eff00;
          16'h13a4 : blkif.rom_rdata <= 32'h938efe0f;
          16'h13a5 : blkif.rom_rdata <= 32'h130e902f;
          16'h13a6 : blkif.rom_rdata <= 32'he31ad10d;
          16'h13a7 : blkif.rom_rdata <= 32'hb7000080;
          16'h13a8 : blkif.rom_rdata <= 32'h93804000;
          16'h13a9 : blkif.rom_rdata <= 32'h1301b02f;
          16'h13aa : blkif.rom_rdata <= 32'h23a02000;
          16'h13ab : blkif.rom_rdata <= 32'hb7101111;
          16'h13ac : blkif.rom_rdata <= 32'h93801011;
          16'h13ad : blkif.rom_rdata <= 32'h37212222;
          16'h13ae : blkif.rom_rdata <= 32'h13012122;
          16'h13af : blkif.rom_rdata <= 32'h33c02000;
          16'h13b0 : blkif.rom_rdata <= 32'h930e0000;
          16'h13b1 : blkif.rom_rdata <= 32'h130eb02f;
          16'h13b2 : blkif.rom_rdata <= 32'he312d00b;
          16'h13b3 : blkif.rom_rdata <= 32'hb7000080;
          16'h13b4 : blkif.rom_rdata <= 32'h93804000;
          16'h13b5 : blkif.rom_rdata <= 32'h1301c02f;
          16'h13b6 : blkif.rom_rdata <= 32'h23a02000;
          16'h13b7 : blkif.rom_rdata <= 32'hb710ff00;
          16'h13b8 : blkif.rom_rdata <= 32'h938000f0;
          16'h13b9 : blkif.rom_rdata <= 32'h93c1f0f0;
          16'h13ba : blkif.rom_rdata <= 32'hb7fe00ff;
          16'h13bb : blkif.rom_rdata <= 32'h938efe00;
          16'h13bc : blkif.rom_rdata <= 32'h130ec02f;
          16'h13bd : blkif.rom_rdata <= 32'he39cd107;
          16'h13be : blkif.rom_rdata <= 32'hb7000080;
          16'h13bf : blkif.rom_rdata <= 32'h93804000;
          16'h13c0 : blkif.rom_rdata <= 32'h1301d02f;
          16'h13c1 : blkif.rom_rdata <= 32'h23a02000;
          16'h13c2 : blkif.rom_rdata <= 32'hb710f00f;
          16'h13c3 : blkif.rom_rdata <= 32'h938000ff;
          16'h13c4 : blkif.rom_rdata <= 32'h93c1000f;
          16'h13c5 : blkif.rom_rdata <= 32'hb71ef00f;
          16'h13c6 : blkif.rom_rdata <= 32'h938e0ef0;
          16'h13c7 : blkif.rom_rdata <= 32'h130ed02f;
          16'h13c8 : blkif.rom_rdata <= 32'he396d105;
          16'h13c9 : blkif.rom_rdata <= 32'hb7000080;
          16'h13ca : blkif.rom_rdata <= 32'h93804000;
          16'h13cb : blkif.rom_rdata <= 32'h13010030;
          16'h13cc : blkif.rom_rdata <= 32'h23a02000;
          16'h13cd : blkif.rom_rdata <= 32'hb7f000ff;
          16'h13ce : blkif.rom_rdata <= 32'h93800070;
          16'h13cf : blkif.rom_rdata <= 32'h93c0f070;
          16'h13d0 : blkif.rom_rdata <= 32'hb7fe00ff;
          16'h13d1 : blkif.rom_rdata <= 32'h938efe00;
          16'h13d2 : blkif.rom_rdata <= 32'h130e0030;
          16'h13d3 : blkif.rom_rdata <= 32'he390d003;
          16'h13d4 : blkif.rom_rdata <= 32'hb7000080;
          16'h13d5 : blkif.rom_rdata <= 32'h93804000;
          16'h13d6 : blkif.rom_rdata <= 32'h13011030;
          16'h13d7 : blkif.rom_rdata <= 32'h23a02000;
          16'h13d8 : blkif.rom_rdata <= 32'h13020000;
          16'h13d9 : blkif.rom_rdata <= 32'hb710f00f;
          16'h13da : blkif.rom_rdata <= 32'h938000ff;
          16'h13db : blkif.rom_rdata <= 32'h93c1000f;
          16'h13dc : blkif.rom_rdata <= 32'h13830100;
          16'h13dd : blkif.rom_rdata <= 32'h13021200;
          16'h13de : blkif.rom_rdata <= 32'h93022000;
          16'h13df : blkif.rom_rdata <= 32'he31452fe;
          16'h13e0 : blkif.rom_rdata <= 32'hb71ef00f;
          16'h13e1 : blkif.rom_rdata <= 32'h938e0ef0;
          16'h13e2 : blkif.rom_rdata <= 32'h130e1030;
          16'h13e3 : blkif.rom_rdata <= 32'h6310d37f;
          16'h13e4 : blkif.rom_rdata <= 32'hb7000080;
          16'h13e5 : blkif.rom_rdata <= 32'h93804000;
          16'h13e6 : blkif.rom_rdata <= 32'h13014030;
          16'h13e7 : blkif.rom_rdata <= 32'h23a02000;
          16'h13e8 : blkif.rom_rdata <= 32'h13020000;
          16'h13e9 : blkif.rom_rdata <= 32'hb710f00f;
          16'h13ea : blkif.rom_rdata <= 32'h938000ff;
          16'h13eb : blkif.rom_rdata <= 32'h93c1000f;
          16'h13ec : blkif.rom_rdata <= 32'h13021200;
          16'h13ed : blkif.rom_rdata <= 32'h93022000;
          16'h13ee : blkif.rom_rdata <= 32'he31652fe;
          16'h13ef : blkif.rom_rdata <= 32'hb71ef00f;
          16'h13f0 : blkif.rom_rdata <= 32'h938e0ef0;
          16'h13f1 : blkif.rom_rdata <= 32'h130e4030;
          16'h13f2 : blkif.rom_rdata <= 32'h6392d17b;
          16'h13f3 : blkif.rom_rdata <= 32'hb7000080;
          16'h13f4 : blkif.rom_rdata <= 32'h93804000;
          16'h13f5 : blkif.rom_rdata <= 32'h13016030;
          16'h13f6 : blkif.rom_rdata <= 32'h23a02000;
          16'h13f7 : blkif.rom_rdata <= 32'h13020000;
          16'h13f8 : blkif.rom_rdata <= 32'hb7f00ff0;
          16'h13f9 : blkif.rom_rdata <= 32'h9380f000;
          16'h13fa : blkif.rom_rdata <= 32'h13000000;
          16'h13fb : blkif.rom_rdata <= 32'h13000000;
          16'h13fc : blkif.rom_rdata <= 32'h93c1000f;
          16'h13fd : blkif.rom_rdata <= 32'h13021200;
          16'h13fe : blkif.rom_rdata <= 32'h93022000;
          16'h13ff : blkif.rom_rdata <= 32'he31252fe;
          16'h1400 : blkif.rom_rdata <= 32'hb7fe0ff0;
          16'h1401 : blkif.rom_rdata <= 32'h938efe0f;
          16'h1402 : blkif.rom_rdata <= 32'h130e6030;
          16'h1403 : blkif.rom_rdata <= 32'h6390d177;
          16'h1404 : blkif.rom_rdata <= 32'hb7000080;
          16'h1405 : blkif.rom_rdata <= 32'h93804000;
          16'h1406 : blkif.rom_rdata <= 32'h13017030;
          16'h1407 : blkif.rom_rdata <= 32'h23a02000;
          16'h1408 : blkif.rom_rdata <= 32'h9340000f;
          16'h1409 : blkif.rom_rdata <= 32'h930e000f;
          16'h140a : blkif.rom_rdata <= 32'h130e7030;
          16'h140b : blkif.rom_rdata <= 32'h6390d075;
          16'h140c : blkif.rom_rdata <= 32'hb7000080;
          16'h140d : blkif.rom_rdata <= 32'h93804000;
          16'h140e : blkif.rom_rdata <= 32'h13018030;
          16'h140f : blkif.rom_rdata <= 32'h23a02000;
          16'h1410 : blkif.rom_rdata <= 32'hb700ff00;
          16'h1411 : blkif.rom_rdata <= 32'h9380f00f;
          16'h1412 : blkif.rom_rdata <= 32'h13c0f070;
          16'h1413 : blkif.rom_rdata <= 32'h930e0000;
          16'h1414 : blkif.rom_rdata <= 32'h130e8030;
          16'h1415 : blkif.rom_rdata <= 32'h631cd071;
          16'h1416 : blkif.rom_rdata <= 32'h130e9030;
          16'h1417 : blkif.rom_rdata <= 32'hb7000080;
          16'h1418 : blkif.rom_rdata <= 32'h93804000;
          16'h1419 : blkif.rom_rdata <= 32'h13019030;
          16'h141a : blkif.rom_rdata <= 32'h23a02000;
          16'h141b : blkif.rom_rdata <= 32'h93610000;
          16'h141c : blkif.rom_rdata <= 32'h13620000;
          16'h141d : blkif.rom_rdata <= 32'h93103000;
          16'h141e : blkif.rom_rdata <= 32'h17110000;
          16'h141f : blkif.rom_rdata <= 32'h130181f8;
          16'h1420 : blkif.rom_rdata <= 32'h33011100;
          16'h1421 : blkif.rom_rdata <= 32'h83200100;
          16'h1422 : blkif.rom_rdata <= 32'h9390e000;
          16'h1423 : blkif.rom_rdata <= 32'h03214100;
          16'h1424 : blkif.rom_rdata <= 32'hb3e02000;
          16'h1425 : blkif.rom_rdata <= 32'h37010090;
          16'h1426 : blkif.rom_rdata <= 32'h23201100;
          16'h1427 : blkif.rom_rdata <= 32'h13000000;
          16'h1428 : blkif.rom_rdata <= 32'h13000000;
          16'h1429 : blkif.rom_rdata <= 32'h13000000;
          16'h142a : blkif.rom_rdata <= 32'h6f00406c;
          16'h142b : blkif.rom_rdata <= 32'h6f00006c;
          16'h142c : blkif.rom_rdata <= 32'h6f00c06b;
          16'h142d : blkif.rom_rdata <= 32'h6f00806b;
          16'h142e : blkif.rom_rdata <= 32'h130ea030;
          16'h142f : blkif.rom_rdata <= 32'hb7000080;
          16'h1430 : blkif.rom_rdata <= 32'h93804000;
          16'h1431 : blkif.rom_rdata <= 32'h1301a030;
          16'h1432 : blkif.rom_rdata <= 32'h23a02000;
          16'h1433 : blkif.rom_rdata <= 32'h93610000;
          16'h1434 : blkif.rom_rdata <= 32'h13620000;
          16'h1435 : blkif.rom_rdata <= 32'h93620000;
          16'h1436 : blkif.rom_rdata <= 32'h9364f001;
          16'h1437 : blkif.rom_rdata <= 32'h17040000;
          16'h1438 : blkif.rom_rdata <= 32'h1304c403;
          16'h1439 : blkif.rom_rdata <= 32'h63c0540e;
          16'h143a : blkif.rom_rdata <= 32'h13933200;
          16'h143b : blkif.rom_rdata <= 32'h97130000;
          16'h143c : blkif.rom_rdata <= 32'h9383c3f1;
          16'h143d : blkif.rom_rdata <= 32'hb3836300;
          16'h143e : blkif.rom_rdata <= 32'h03a30300;
          16'h143f : blkif.rom_rdata <= 32'h1313e300;
          16'h1440 : blkif.rom_rdata <= 32'h83a34300;
          16'h1441 : blkif.rom_rdata <= 32'h33637300;
          16'h1442 : blkif.rom_rdata <= 32'hb7030090;
          16'h1443 : blkif.rom_rdata <= 32'h23a06300;
          16'h1444 : blkif.rom_rdata <= 32'h13000000;
          16'h1445 : blkif.rom_rdata <= 32'h13000000;
          16'h1446 : blkif.rom_rdata <= 32'h13000000;
          16'h1447 : blkif.rom_rdata <= 32'hef004009;
          16'h1448 : blkif.rom_rdata <= 32'hef000009;
          16'h1449 : blkif.rom_rdata <= 32'hef00c008;
          16'h144a : blkif.rom_rdata <= 32'hef008008;
          16'h144b : blkif.rom_rdata <= 32'hef004008;
          16'h144c : blkif.rom_rdata <= 32'hef000008;
          16'h144d : blkif.rom_rdata <= 32'hef00c007;
          16'h144e : blkif.rom_rdata <= 32'hef008007;
          16'h144f : blkif.rom_rdata <= 32'hef004007;
          16'h1450 : blkif.rom_rdata <= 32'hef000007;
          16'h1451 : blkif.rom_rdata <= 32'hef00c006;
          16'h1452 : blkif.rom_rdata <= 32'hef008006;
          16'h1453 : blkif.rom_rdata <= 32'hef004006;
          16'h1454 : blkif.rom_rdata <= 32'hef000006;
          16'h1455 : blkif.rom_rdata <= 32'hef00c005;
          16'h1456 : blkif.rom_rdata <= 32'hef008005;
          16'h1457 : blkif.rom_rdata <= 32'hef004005;
          16'h1458 : blkif.rom_rdata <= 32'hef000005;
          16'h1459 : blkif.rom_rdata <= 32'hef00c004;
          16'h145a : blkif.rom_rdata <= 32'hef008004;
          16'h145b : blkif.rom_rdata <= 32'hef004004;
          16'h145c : blkif.rom_rdata <= 32'hef000004;
          16'h145d : blkif.rom_rdata <= 32'hef00c003;
          16'h145e : blkif.rom_rdata <= 32'hef008003;
          16'h145f : blkif.rom_rdata <= 32'hef004003;
          16'h1460 : blkif.rom_rdata <= 32'hef000003;
          16'h1461 : blkif.rom_rdata <= 32'hef00c002;
          16'h1462 : blkif.rom_rdata <= 32'hef008002;
          16'h1463 : blkif.rom_rdata <= 32'hef004002;
          16'h1464 : blkif.rom_rdata <= 32'hef000002;
          16'h1465 : blkif.rom_rdata <= 32'hef00c001;
          16'h1466 : blkif.rom_rdata <= 32'hef008001;
          16'h1467 : blkif.rom_rdata <= 32'h6f00005d;
          16'h1468 : blkif.rom_rdata <= 32'h6f00c05c;
          16'h1469 : blkif.rom_rdata <= 32'h6f00805c;
          16'h146a : blkif.rom_rdata <= 32'h6f00405c;
          16'h146b : blkif.rom_rdata <= 32'h6f00005c;
          16'h146c : blkif.rom_rdata <= 32'h13952200;
          16'h146d : blkif.rom_rdata <= 32'h938080ff;
          16'h146e : blkif.rom_rdata <= 32'hb380a040;
          16'h146f : blkif.rom_rdata <= 32'h93821200;
          16'h1470 : blkif.rom_rdata <= 32'he38280f2;
          16'h1471 : blkif.rom_rdata <= 32'h130eb030;
          16'h1472 : blkif.rom_rdata <= 32'hb7000080;
          16'h1473 : blkif.rom_rdata <= 32'h93804000;
          16'h1474 : blkif.rom_rdata <= 32'h1301b030;
          16'h1475 : blkif.rom_rdata <= 32'h23a02000;
          16'h1476 : blkif.rom_rdata <= 32'h93611000;
          16'h1477 : blkif.rom_rdata <= 32'h13620000;
          16'h1478 : blkif.rom_rdata <= 32'h93620000;
          16'h1479 : blkif.rom_rdata <= 32'h13933200;
          16'h147a : blkif.rom_rdata <= 32'h97130000;
          16'h147b : blkif.rom_rdata <= 32'h938303f2;
          16'h147c : blkif.rom_rdata <= 32'hb3836300;
          16'h147d : blkif.rom_rdata <= 32'h03a30300;
          16'h147e : blkif.rom_rdata <= 32'h1313e300;
          16'h147f : blkif.rom_rdata <= 32'h83a34300;
          16'h1480 : blkif.rom_rdata <= 32'h33637300;
          16'h1481 : blkif.rom_rdata <= 32'hb7030090;
          16'h1482 : blkif.rom_rdata <= 32'h23a06300;
          16'h1483 : blkif.rom_rdata <= 32'h93821200;
          16'h1484 : blkif.rom_rdata <= 32'h13933200;
          16'h1485 : blkif.rom_rdata <= 32'h97130000;
          16'h1486 : blkif.rom_rdata <= 32'h938343ef;
          16'h1487 : blkif.rom_rdata <= 32'hb3836300;
          16'h1488 : blkif.rom_rdata <= 32'h03a30300;
          16'h1489 : blkif.rom_rdata <= 32'h1313e300;
          16'h148a : blkif.rom_rdata <= 32'h83a34300;
          16'h148b : blkif.rom_rdata <= 32'h33637300;
          16'h148c : blkif.rom_rdata <= 32'hb7030090;
          16'h148d : blkif.rom_rdata <= 32'h23a06300;
          16'h148e : blkif.rom_rdata <= 32'h93821200;
          16'h148f : blkif.rom_rdata <= 32'h13933200;
          16'h1490 : blkif.rom_rdata <= 32'h97130000;
          16'h1491 : blkif.rom_rdata <= 32'h938383ec;
          16'h1492 : blkif.rom_rdata <= 32'hb3836300;
          16'h1493 : blkif.rom_rdata <= 32'h03a30300;
          16'h1494 : blkif.rom_rdata <= 32'h1313e300;
          16'h1495 : blkif.rom_rdata <= 32'h83a34300;
          16'h1496 : blkif.rom_rdata <= 32'h33637300;
          16'h1497 : blkif.rom_rdata <= 32'hb7030090;
          16'h1498 : blkif.rom_rdata <= 32'h23a06300;
          16'h1499 : blkif.rom_rdata <= 32'h93821200;
          16'h149a : blkif.rom_rdata <= 32'h13933200;
          16'h149b : blkif.rom_rdata <= 32'h97130000;
          16'h149c : blkif.rom_rdata <= 32'h9383c3e9;
          16'h149d : blkif.rom_rdata <= 32'hb3836300;
          16'h149e : blkif.rom_rdata <= 32'h03a30300;
          16'h149f : blkif.rom_rdata <= 32'h1313e300;
          16'h14a0 : blkif.rom_rdata <= 32'h83a34300;
          16'h14a1 : blkif.rom_rdata <= 32'h33637300;
          16'h14a2 : blkif.rom_rdata <= 32'hb7030090;
          16'h14a3 : blkif.rom_rdata <= 32'h23a06300;
          16'h14a4 : blkif.rom_rdata <= 32'h13000000;
          16'h14a5 : blkif.rom_rdata <= 32'h13000000;
          16'h14a6 : blkif.rom_rdata <= 32'h93610000;
          16'h14a7 : blkif.rom_rdata <= 32'h13000000;
          16'h14a8 : blkif.rom_rdata <= 32'h6f00c04c;
          16'h14a9 : blkif.rom_rdata <= 32'h6f00804c;
          16'h14aa : blkif.rom_rdata <= 32'h6312304c;
          16'h14ab : blkif.rom_rdata <= 32'h13621000;
          16'h14ac : blkif.rom_rdata <= 32'h63164000;
          16'h14ad : blkif.rom_rdata <= 32'h6f00804b;
          16'h14ae : blkif.rom_rdata <= 32'h6f00404b;
          16'h14af : blkif.rom_rdata <= 32'h93611000;
          16'h14b0 : blkif.rom_rdata <= 32'h63164000;
          16'h14b1 : blkif.rom_rdata <= 32'h6f00804a;
          16'h14b2 : blkif.rom_rdata <= 32'h6f00404a;
          16'h14b3 : blkif.rom_rdata <= 32'h93610000;
          16'h14b4 : blkif.rom_rdata <= 32'h13000000;
          16'h14b5 : blkif.rom_rdata <= 32'h6f008049;
          16'h14b6 : blkif.rom_rdata <= 32'h6f004049;
          16'h14b7 : blkif.rom_rdata <= 32'h130ec030;
          16'h14b8 : blkif.rom_rdata <= 32'hb7000080;
          16'h14b9 : blkif.rom_rdata <= 32'h93804000;
          16'h14ba : blkif.rom_rdata <= 32'h1301c030;
          16'h14bb : blkif.rom_rdata <= 32'h23a02000;
          16'h14bc : blkif.rom_rdata <= 32'h93610000;
          16'h14bd : blkif.rom_rdata <= 32'h13620000;
          16'h14be : blkif.rom_rdata <= 32'h93620000;
          16'h14bf : blkif.rom_rdata <= 32'h13933200;
          16'h14c0 : blkif.rom_rdata <= 32'h97130000;
          16'h14c1 : blkif.rom_rdata <= 32'h938383e2;
          16'h14c2 : blkif.rom_rdata <= 32'hb3836300;
          16'h14c3 : blkif.rom_rdata <= 32'h03a30300;
          16'h14c4 : blkif.rom_rdata <= 32'h1313e300;
          16'h14c5 : blkif.rom_rdata <= 32'h83a34300;
          16'h14c6 : blkif.rom_rdata <= 32'h33637300;
          16'h14c7 : blkif.rom_rdata <= 32'hb7030090;
          16'h14c8 : blkif.rom_rdata <= 32'h23a06300;
          16'h14c9 : blkif.rom_rdata <= 32'h93821200;
          16'h14ca : blkif.rom_rdata <= 32'h13933200;
          16'h14cb : blkif.rom_rdata <= 32'h97130000;
          16'h14cc : blkif.rom_rdata <= 32'h9383c3df;
          16'h14cd : blkif.rom_rdata <= 32'hb3836300;
          16'h14ce : blkif.rom_rdata <= 32'h03a30300;
          16'h14cf : blkif.rom_rdata <= 32'h1313e300;
          16'h14d0 : blkif.rom_rdata <= 32'h83a34300;
          16'h14d1 : blkif.rom_rdata <= 32'h33637300;
          16'h14d2 : blkif.rom_rdata <= 32'hb7030090;
          16'h14d3 : blkif.rom_rdata <= 32'h23a06300;
          16'h14d4 : blkif.rom_rdata <= 32'h93821200;
          16'h14d5 : blkif.rom_rdata <= 32'h13933200;
          16'h14d6 : blkif.rom_rdata <= 32'h97130000;
          16'h14d7 : blkif.rom_rdata <= 32'h938303dd;
          16'h14d8 : blkif.rom_rdata <= 32'hb3836300;
          16'h14d9 : blkif.rom_rdata <= 32'h03a30300;
          16'h14da : blkif.rom_rdata <= 32'h1313e300;
          16'h14db : blkif.rom_rdata <= 32'h83a34300;
          16'h14dc : blkif.rom_rdata <= 32'h33637300;
          16'h14dd : blkif.rom_rdata <= 32'hb7030090;
          16'h14de : blkif.rom_rdata <= 32'h23a06300;
          16'h14df : blkif.rom_rdata <= 32'h93821200;
          16'h14e0 : blkif.rom_rdata <= 32'h13933200;
          16'h14e1 : blkif.rom_rdata <= 32'h97130000;
          16'h14e2 : blkif.rom_rdata <= 32'h938343da;
          16'h14e3 : blkif.rom_rdata <= 32'hb3836300;
          16'h14e4 : blkif.rom_rdata <= 32'h03a30300;
          16'h14e5 : blkif.rom_rdata <= 32'h1313e300;
          16'h14e6 : blkif.rom_rdata <= 32'h83a34300;
          16'h14e7 : blkif.rom_rdata <= 32'h33637300;
          16'h14e8 : blkif.rom_rdata <= 32'hb7030090;
          16'h14e9 : blkif.rom_rdata <= 32'h23a06300;
          16'h14ea : blkif.rom_rdata <= 32'h13000000;
          16'h14eb : blkif.rom_rdata <= 32'h13000000;
          16'h14ec : blkif.rom_rdata <= 32'h93611000;
          16'h14ed : blkif.rom_rdata <= 32'h6f00803b;
          16'h14ee : blkif.rom_rdata <= 32'h6f00403b;
          16'h14ef : blkif.rom_rdata <= 32'h6308303a;
          16'h14f0 : blkif.rom_rdata <= 32'h93610000;
          16'h14f1 : blkif.rom_rdata <= 32'h63083000;
          16'h14f2 : blkif.rom_rdata <= 32'h6f00403a;
          16'h14f3 : blkif.rom_rdata <= 32'h6f00003a;
          16'h14f4 : blkif.rom_rdata <= 32'h6f00c039;
          16'h14f5 : blkif.rom_rdata <= 32'h93611000;
          16'h14f6 : blkif.rom_rdata <= 32'h6f004039;
          16'h14f7 : blkif.rom_rdata <= 32'h6f000039;
          16'h14f8 : blkif.rom_rdata <= 32'h13621000;
          16'h14f9 : blkif.rom_rdata <= 32'h63043038;
          16'h14fa : blkif.rom_rdata <= 32'h93610000;
          16'h14fb : blkif.rom_rdata <= 32'h63083000;
          16'h14fc : blkif.rom_rdata <= 32'h6f00c037;
          16'h14fd : blkif.rom_rdata <= 32'h6f008037;
          16'h14fe : blkif.rom_rdata <= 32'h6f004037;
          16'h14ff : blkif.rom_rdata <= 32'h130ed030;
          16'h1500 : blkif.rom_rdata <= 32'hb7000080;
          16'h1501 : blkif.rom_rdata <= 32'h93804000;
          16'h1502 : blkif.rom_rdata <= 32'h1301d030;
          16'h1503 : blkif.rom_rdata <= 32'h23a02000;
          16'h1504 : blkif.rom_rdata <= 32'h93610000;
          16'h1505 : blkif.rom_rdata <= 32'h13620000;
          16'h1506 : blkif.rom_rdata <= 32'h93620000;
          16'h1507 : blkif.rom_rdata <= 32'h13933200;
          16'h1508 : blkif.rom_rdata <= 32'h97130000;
          16'h1509 : blkif.rom_rdata <= 32'h938383d2;
          16'h150a : blkif.rom_rdata <= 32'hb3836300;
          16'h150b : blkif.rom_rdata <= 32'h03a30300;
          16'h150c : blkif.rom_rdata <= 32'h1313e300;
          16'h150d : blkif.rom_rdata <= 32'h83a34300;
          16'h150e : blkif.rom_rdata <= 32'h33637300;
          16'h150f : blkif.rom_rdata <= 32'hb7030090;
          16'h1510 : blkif.rom_rdata <= 32'h23a06300;
          16'h1511 : blkif.rom_rdata <= 32'h93821200;
          16'h1512 : blkif.rom_rdata <= 32'h13933200;
          16'h1513 : blkif.rom_rdata <= 32'h97130000;
          16'h1514 : blkif.rom_rdata <= 32'h9383c3cf;
          16'h1515 : blkif.rom_rdata <= 32'hb3836300;
          16'h1516 : blkif.rom_rdata <= 32'h03a30300;
          16'h1517 : blkif.rom_rdata <= 32'h1313e300;
          16'h1518 : blkif.rom_rdata <= 32'h83a34300;
          16'h1519 : blkif.rom_rdata <= 32'h33637300;
          16'h151a : blkif.rom_rdata <= 32'hb7030090;
          16'h151b : blkif.rom_rdata <= 32'h23a06300;
          16'h151c : blkif.rom_rdata <= 32'h93821200;
          16'h151d : blkif.rom_rdata <= 32'h13933200;
          16'h151e : blkif.rom_rdata <= 32'h97130000;
          16'h151f : blkif.rom_rdata <= 32'h938303cd;
          16'h1520 : blkif.rom_rdata <= 32'hb3836300;
          16'h1521 : blkif.rom_rdata <= 32'h03a30300;
          16'h1522 : blkif.rom_rdata <= 32'h1313e300;
          16'h1523 : blkif.rom_rdata <= 32'h83a34300;
          16'h1524 : blkif.rom_rdata <= 32'h33637300;
          16'h1525 : blkif.rom_rdata <= 32'hb7030090;
          16'h1526 : blkif.rom_rdata <= 32'h23a06300;
          16'h1527 : blkif.rom_rdata <= 32'h93821200;
          16'h1528 : blkif.rom_rdata <= 32'h13933200;
          16'h1529 : blkif.rom_rdata <= 32'h97130000;
          16'h152a : blkif.rom_rdata <= 32'h938343ca;
          16'h152b : blkif.rom_rdata <= 32'hb3836300;
          16'h152c : blkif.rom_rdata <= 32'h03a30300;
          16'h152d : blkif.rom_rdata <= 32'h1313e300;
          16'h152e : blkif.rom_rdata <= 32'h83a34300;
          16'h152f : blkif.rom_rdata <= 32'h33637300;
          16'h1530 : blkif.rom_rdata <= 32'hb7030090;
          16'h1531 : blkif.rom_rdata <= 32'h23a06300;
          16'h1532 : blkif.rom_rdata <= 32'h93821200;
          16'h1533 : blkif.rom_rdata <= 32'h13933200;
          16'h1534 : blkif.rom_rdata <= 32'h97130000;
          16'h1535 : blkif.rom_rdata <= 32'h938383c7;
          16'h1536 : blkif.rom_rdata <= 32'hb3836300;
          16'h1537 : blkif.rom_rdata <= 32'h03a30300;
          16'h1538 : blkif.rom_rdata <= 32'h1313e300;
          16'h1539 : blkif.rom_rdata <= 32'h83a34300;
          16'h153a : blkif.rom_rdata <= 32'h33637300;
          16'h153b : blkif.rom_rdata <= 32'hb7030090;
          16'h153c : blkif.rom_rdata <= 32'h23a06300;
          16'h153d : blkif.rom_rdata <= 32'h13000000;
          16'h153e : blkif.rom_rdata <= 32'h13000000;
          16'h153f : blkif.rom_rdata <= 32'h97020000;
          16'h1540 : blkif.rom_rdata <= 32'h9382c202;
          16'h1541 : blkif.rom_rdata <= 32'h13647000;
          16'h1542 : blkif.rom_rdata <= 32'h6f00c000;
          16'h1543 : blkif.rom_rdata <= 32'h6f000026;
          16'h1544 : blkif.rom_rdata <= 32'h6f00c025;
          16'h1545 : blkif.rom_rdata <= 32'he7800200;
          16'h1546 : blkif.rom_rdata <= 32'h6f004025;
          16'h1547 : blkif.rom_rdata <= 32'h6f000025;
          16'h1548 : blkif.rom_rdata <= 32'h6f00c024;
          16'h1549 : blkif.rom_rdata <= 32'h6f008024;
          16'h154a : blkif.rom_rdata <= 32'h63060000;
          16'h154b : blkif.rom_rdata <= 32'h6f000024;
          16'h154c : blkif.rom_rdata <= 32'h6f00c023;
          16'h154d : blkif.rom_rdata <= 32'h631a8000;
          16'h154e : blkif.rom_rdata <= 32'h6f004023;
          16'h154f : blkif.rom_rdata <= 32'h6f000023;
          16'h1550 : blkif.rom_rdata <= 32'h6f00c022;
          16'h1551 : blkif.rom_rdata <= 32'h6f008022;
          16'h1552 : blkif.rom_rdata <= 32'h63468000;
          16'h1553 : blkif.rom_rdata <= 32'h6f000022;
          16'h1554 : blkif.rom_rdata <= 32'h6f00c021;
          16'h1555 : blkif.rom_rdata <= 32'h130ee030;
          16'h1556 : blkif.rom_rdata <= 32'hb7000080;
          16'h1557 : blkif.rom_rdata <= 32'h93804000;
          16'h1558 : blkif.rom_rdata <= 32'h1301e030;
          16'h1559 : blkif.rom_rdata <= 32'h23a02000;
          16'h155a : blkif.rom_rdata <= 32'h93610000;
          16'h155b : blkif.rom_rdata <= 32'h13620000;
          16'h155c : blkif.rom_rdata <= 32'h93620000;
          16'h155d : blkif.rom_rdata <= 32'h13933200;
          16'h155e : blkif.rom_rdata <= 32'h97130000;
          16'h155f : blkif.rom_rdata <= 32'h938383bf;
          16'h1560 : blkif.rom_rdata <= 32'hb3836300;
          16'h1561 : blkif.rom_rdata <= 32'h03a30300;
          16'h1562 : blkif.rom_rdata <= 32'h1313e300;
          16'h1563 : blkif.rom_rdata <= 32'h83a34300;
          16'h1564 : blkif.rom_rdata <= 32'h33637300;
          16'h1565 : blkif.rom_rdata <= 32'hb7030090;
          16'h1566 : blkif.rom_rdata <= 32'h23a06300;
          16'h1567 : blkif.rom_rdata <= 32'h93821200;
          16'h1568 : blkif.rom_rdata <= 32'h13933200;
          16'h1569 : blkif.rom_rdata <= 32'h97130000;
          16'h156a : blkif.rom_rdata <= 32'h9383c3bc;
          16'h156b : blkif.rom_rdata <= 32'hb3836300;
          16'h156c : blkif.rom_rdata <= 32'h03a30300;
          16'h156d : blkif.rom_rdata <= 32'h1313e300;
          16'h156e : blkif.rom_rdata <= 32'h83a34300;
          16'h156f : blkif.rom_rdata <= 32'h33637300;
          16'h1570 : blkif.rom_rdata <= 32'hb7030090;
          16'h1571 : blkif.rom_rdata <= 32'h23a06300;
          16'h1572 : blkif.rom_rdata <= 32'h93821200;
          16'h1573 : blkif.rom_rdata <= 32'h13933200;
          16'h1574 : blkif.rom_rdata <= 32'h97130000;
          16'h1575 : blkif.rom_rdata <= 32'h938303ba;
          16'h1576 : blkif.rom_rdata <= 32'hb3836300;
          16'h1577 : blkif.rom_rdata <= 32'h03a30300;
          16'h1578 : blkif.rom_rdata <= 32'h1313e300;
          16'h1579 : blkif.rom_rdata <= 32'h83a34300;
          16'h157a : blkif.rom_rdata <= 32'h33637300;
          16'h157b : blkif.rom_rdata <= 32'hb7030090;
          16'h157c : blkif.rom_rdata <= 32'h23a06300;
          16'h157d : blkif.rom_rdata <= 32'h13000000;
          16'h157e : blkif.rom_rdata <= 32'h13000000;
          16'h157f : blkif.rom_rdata <= 32'h63180016;
          16'h1580 : blkif.rom_rdata <= 32'h6f008000;
          16'h1581 : blkif.rom_rdata <= 32'h6f008016;
          16'h1582 : blkif.rom_rdata <= 32'h63820216;
          16'h1583 : blkif.rom_rdata <= 32'h6f000001;
          16'h1584 : blkif.rom_rdata <= 32'h6f00c015;
          16'h1585 : blkif.rom_rdata <= 32'h6f008015;
          16'h1586 : blkif.rom_rdata <= 32'h6f004015;
          16'h1587 : blkif.rom_rdata <= 32'h63c80214;
          16'h1588 : blkif.rom_rdata <= 32'h6f008000;
          16'h1589 : blkif.rom_rdata <= 32'h6f008014;
          16'h158a : blkif.rom_rdata <= 32'h130ef030;
          16'h158b : blkif.rom_rdata <= 32'hb7000080;
          16'h158c : blkif.rom_rdata <= 32'h93804000;
          16'h158d : blkif.rom_rdata <= 32'h1301f030;
          16'h158e : blkif.rom_rdata <= 32'h23a02000;
          16'h158f : blkif.rom_rdata <= 32'h93610000;
          16'h1590 : blkif.rom_rdata <= 32'h13620000;
          16'h1591 : blkif.rom_rdata <= 32'h93620000;
          16'h1592 : blkif.rom_rdata <= 32'h13933200;
          16'h1593 : blkif.rom_rdata <= 32'h97130000;
          16'h1594 : blkif.rom_rdata <= 32'h9383c3b3;
          16'h1595 : blkif.rom_rdata <= 32'hb3836300;
          16'h1596 : blkif.rom_rdata <= 32'h03a30300;
          16'h1597 : blkif.rom_rdata <= 32'h1313e300;
          16'h1598 : blkif.rom_rdata <= 32'h83a34300;
          16'h1599 : blkif.rom_rdata <= 32'h33637300;
          16'h159a : blkif.rom_rdata <= 32'hb7030090;
          16'h159b : blkif.rom_rdata <= 32'h23a06300;
          16'h159c : blkif.rom_rdata <= 32'h93821200;
          16'h159d : blkif.rom_rdata <= 32'h13000000;
          16'h159e : blkif.rom_rdata <= 32'h13000000;
          16'h159f : blkif.rom_rdata <= 32'h13000000;
          16'h15a0 : blkif.rom_rdata <= 32'h13000000;
          16'h15a1 : blkif.rom_rdata <= 32'h6f00800e;
          16'h15a2 : blkif.rom_rdata <= 32'h6f00400e;
          16'h15a3 : blkif.rom_rdata <= 32'h37040090;
          16'h15a4 : blkif.rom_rdata <= 32'h13044400;
          16'h15a5 : blkif.rom_rdata <= 32'h23205400;
          16'h15a6 : blkif.rom_rdata <= 32'h13933200;
          16'h15a7 : blkif.rom_rdata <= 32'h97130000;
          16'h15a8 : blkif.rom_rdata <= 32'h9383c3ae;
          16'h15a9 : blkif.rom_rdata <= 32'hb3836300;
          16'h15aa : blkif.rom_rdata <= 32'h03a30300;
          16'h15ab : blkif.rom_rdata <= 32'h1313e300;
          16'h15ac : blkif.rom_rdata <= 32'h83a34300;
          16'h15ad : blkif.rom_rdata <= 32'h33637300;
          16'h15ae : blkif.rom_rdata <= 32'hb7030090;
          16'h15af : blkif.rom_rdata <= 32'h23a06300;
          16'h15b0 : blkif.rom_rdata <= 32'h93821200;
          16'h15b1 : blkif.rom_rdata <= 32'h13933200;
          16'h15b2 : blkif.rom_rdata <= 32'h97130000;
          16'h15b3 : blkif.rom_rdata <= 32'h938303ac;
          16'h15b4 : blkif.rom_rdata <= 32'hb3836300;
          16'h15b5 : blkif.rom_rdata <= 32'h03a30300;
          16'h15b6 : blkif.rom_rdata <= 32'h1313e300;
          16'h15b7 : blkif.rom_rdata <= 32'h83a34300;
          16'h15b8 : blkif.rom_rdata <= 32'h33637300;
          16'h15b9 : blkif.rom_rdata <= 32'hb7030090;
          16'h15ba : blkif.rom_rdata <= 32'h23a06300;
          16'h15bb : blkif.rom_rdata <= 32'h93821200;
          16'h15bc : blkif.rom_rdata <= 32'h13933200;
          16'h15bd : blkif.rom_rdata <= 32'h97130000;
          16'h15be : blkif.rom_rdata <= 32'h938343a9;
          16'h15bf : blkif.rom_rdata <= 32'hb3836300;
          16'h15c0 : blkif.rom_rdata <= 32'h03a30300;
          16'h15c1 : blkif.rom_rdata <= 32'h1313e300;
          16'h15c2 : blkif.rom_rdata <= 32'h83a34300;
          16'h15c3 : blkif.rom_rdata <= 32'h33637300;
          16'h15c4 : blkif.rom_rdata <= 32'hb7030090;
          16'h15c5 : blkif.rom_rdata <= 32'h23a06300;
          16'h15c6 : blkif.rom_rdata <= 32'h13000000;
          16'h15c7 : blkif.rom_rdata <= 32'h6f004001;
          16'h15c8 : blkif.rom_rdata <= 32'h6f00c004;
          16'h15c9 : blkif.rom_rdata <= 32'h6f008004;
          16'h15ca : blkif.rom_rdata <= 32'h6f004004;
          16'h15cb : blkif.rom_rdata <= 32'h6f000004;
          16'h15cc : blkif.rom_rdata <= 32'h13000000;
          16'h15cd : blkif.rom_rdata <= 32'h23200400;
          16'h15ce : blkif.rom_rdata <= 32'h6f004001;
          16'h15cf : blkif.rom_rdata <= 32'h6f000003;
          16'h15d0 : blkif.rom_rdata <= 32'h6f00c002;
          16'h15d1 : blkif.rom_rdata <= 32'h6f008002;
          16'h15d2 : blkif.rom_rdata <= 32'h6f004002;
          16'h15d3 : blkif.rom_rdata <= 32'h13000000;
          16'h15d4 : blkif.rom_rdata <= 32'h6f00c001;
          16'h15d5 : blkif.rom_rdata <= 32'h6f008001;
          16'h15d6 : blkif.rom_rdata <= 32'hb7000080;
          16'h15d7 : blkif.rom_rdata <= 32'h93804000;
          16'h15d8 : blkif.rom_rdata <= 32'h1301a00a;
          16'h15d9 : blkif.rom_rdata <= 32'h23a02000;
          16'h15da : blkif.rom_rdata <= 32'h631cc001;
          16'h15db : blkif.rom_rdata <= 32'h0f00f00f;
          16'h15dc : blkif.rom_rdata <= 32'h63000e00;
          16'h15dd : blkif.rom_rdata <= 32'h131e1e00;
          16'h15de : blkif.rom_rdata <= 32'h136e1e00;
          16'h15df : blkif.rom_rdata <= 32'h6f000002;
          16'h15e0 : blkif.rom_rdata <= 32'h0f00f00f;
          16'h15e1 : blkif.rom_rdata <= 32'h130e1000;
          16'h15e2 : blkif.rom_rdata <= 32'h6f004001;
          16'h15e3 : blkif.rom_rdata <= 32'h93001000;
          16'h15e4 : blkif.rom_rdata <= 32'h13011000;
          16'h15e5 : blkif.rom_rdata <= 32'h97300000;
          16'h15e6 : blkif.rom_rdata <= 32'h23a6208e;
          16'h15e7 : blkif.rom_rdata <= 32'h6fa05fa6;
          16'h15e8 : blkif.rom_rdata <= 32'h00000000;
          16'h15e9 : blkif.rom_rdata <= 32'h00000000;
          16'h15ea : blkif.rom_rdata <= 32'h00000000;
          16'h15eb : blkif.rom_rdata <= 32'h00000000;
          16'h15ec : blkif.rom_rdata <= 32'h00000000;
          16'h15ed : blkif.rom_rdata <= 32'h00000000;
          16'h15ee : blkif.rom_rdata <= 32'h00000000;
          16'h15ef : blkif.rom_rdata <= 32'h00000000;
          16'h15f0 : blkif.rom_rdata <= 32'h00000000;
          16'h15f1 : blkif.rom_rdata <= 32'h00000000;
          16'h15f2 : blkif.rom_rdata <= 32'h00000000;
          16'h15f3 : blkif.rom_rdata <= 32'h00000000;
          16'h15f4 : blkif.rom_rdata <= 32'h00000000;
          16'h15f5 : blkif.rom_rdata <= 32'h00000000;
          16'h15f6 : blkif.rom_rdata <= 32'h00000000;
          16'h15f7 : blkif.rom_rdata <= 32'h00000000;
          16'h15f8 : blkif.rom_rdata <= 32'h00000000;
          16'h15f9 : blkif.rom_rdata <= 32'h00000000;
          16'h15fa : blkif.rom_rdata <= 32'h00000000;
          16'h15fb : blkif.rom_rdata <= 32'h00000000;
          16'h15fc : blkif.rom_rdata <= 32'h00000000;
          16'h15fd : blkif.rom_rdata <= 32'h00000000;
          16'h15fe : blkif.rom_rdata <= 32'h00000000;
          16'h15ff : blkif.rom_rdata <= 32'h00000000;
          16'h1600 : blkif.rom_rdata <= 32'h00000000;
          16'h1601 : blkif.rom_rdata <= 32'h00000000;
          16'h1602 : blkif.rom_rdata <= 32'h00000000;
          16'h1603 : blkif.rom_rdata <= 32'h00000000;
          16'h1604 : blkif.rom_rdata <= 32'h00000000;
          16'h1605 : blkif.rom_rdata <= 32'h00000000;
          16'h1606 : blkif.rom_rdata <= 32'h00000000;
          16'h1607 : blkif.rom_rdata <= 32'h00000000;
          16'h1608 : blkif.rom_rdata <= 32'h00000000;
          16'h1609 : blkif.rom_rdata <= 32'h00000000;
          16'h160a : blkif.rom_rdata <= 32'h00000000;
          16'h160b : blkif.rom_rdata <= 32'h00000000;
          16'h160c : blkif.rom_rdata <= 32'h00000000;
          16'h160d : blkif.rom_rdata <= 32'h00000000;
          16'h160e : blkif.rom_rdata <= 32'h00000000;
          16'h160f : blkif.rom_rdata <= 32'h00000000;
          16'h1610 : blkif.rom_rdata <= 32'h00000000;
          16'h1611 : blkif.rom_rdata <= 32'h00000000;
          16'h1612 : blkif.rom_rdata <= 32'h00000000;
          16'h1613 : blkif.rom_rdata <= 32'h00000000;
          16'h1614 : blkif.rom_rdata <= 32'h00000000;
          16'h1615 : blkif.rom_rdata <= 32'h00000000;
          16'h1616 : blkif.rom_rdata <= 32'h00000000;
          16'h1617 : blkif.rom_rdata <= 32'h00000000;
          16'h1618 : blkif.rom_rdata <= 32'h00000000;
          16'h1619 : blkif.rom_rdata <= 32'h00000000;
          16'h161a : blkif.rom_rdata <= 32'h00000000;
          16'h161b : blkif.rom_rdata <= 32'h00000000;
          16'h161c : blkif.rom_rdata <= 32'h00000000;
          16'h161d : blkif.rom_rdata <= 32'h00000000;
          16'h161e : blkif.rom_rdata <= 32'h00000000;
          16'h161f : blkif.rom_rdata <= 32'h00000000;
          16'h1620 : blkif.rom_rdata <= 32'h00000000;
          16'h1621 : blkif.rom_rdata <= 32'h00000000;
          16'h1622 : blkif.rom_rdata <= 32'h00000000;
          16'h1623 : blkif.rom_rdata <= 32'h00000000;
          16'h1624 : blkif.rom_rdata <= 32'h00000000;
          16'h1625 : blkif.rom_rdata <= 32'h00000000;
          16'h1626 : blkif.rom_rdata <= 32'h00000000;
          16'h1627 : blkif.rom_rdata <= 32'h00000000;
          16'h1628 : blkif.rom_rdata <= 32'h00000000;
          16'h1629 : blkif.rom_rdata <= 32'h00000000;
          16'h162a : blkif.rom_rdata <= 32'h00000000;
          16'h162b : blkif.rom_rdata <= 32'h00000000;
          16'h162c : blkif.rom_rdata <= 32'h00000000;
          16'h162d : blkif.rom_rdata <= 32'h00000000;
          16'h162e : blkif.rom_rdata <= 32'h00000000;
          16'h162f : blkif.rom_rdata <= 32'h00000000;
          16'h1630 : blkif.rom_rdata <= 32'h00000000;
          16'h1631 : blkif.rom_rdata <= 32'h00000000;
          16'h1632 : blkif.rom_rdata <= 32'h00000000;
          16'h1633 : blkif.rom_rdata <= 32'h00000000;
          16'h1634 : blkif.rom_rdata <= 32'h00000000;
          16'h1635 : blkif.rom_rdata <= 32'h00000000;
          16'h1636 : blkif.rom_rdata <= 32'h00000000;
          16'h1637 : blkif.rom_rdata <= 32'h00000000;
          16'h1638 : blkif.rom_rdata <= 32'h00000000;
          16'h1639 : blkif.rom_rdata <= 32'h00000000;
          16'h163a : blkif.rom_rdata <= 32'h00000000;
          16'h163b : blkif.rom_rdata <= 32'h00000000;
          16'h163c : blkif.rom_rdata <= 32'h00000000;
          16'h163d : blkif.rom_rdata <= 32'h00000000;
          16'h163e : blkif.rom_rdata <= 32'h00000000;
          16'h163f : blkif.rom_rdata <= 32'h00000000;
          16'h1640 : blkif.rom_rdata <= 32'h00000000;
          16'h1641 : blkif.rom_rdata <= 32'h00000000;
          16'h1642 : blkif.rom_rdata <= 32'h00000000;
          16'h1643 : blkif.rom_rdata <= 32'h00000000;
          16'h1644 : blkif.rom_rdata <= 32'h00000000;
          16'h1645 : blkif.rom_rdata <= 32'h00000000;
          16'h1646 : blkif.rom_rdata <= 32'h00000000;
          16'h1647 : blkif.rom_rdata <= 32'h00000000;
          16'h1648 : blkif.rom_rdata <= 32'h00000000;
          16'h1649 : blkif.rom_rdata <= 32'h00000000;
          16'h164a : blkif.rom_rdata <= 32'h00000000;
          16'h164b : blkif.rom_rdata <= 32'h00000000;
          16'h164c : blkif.rom_rdata <= 32'h00000000;
          16'h164d : blkif.rom_rdata <= 32'h00000000;
          16'h164e : blkif.rom_rdata <= 32'h00000000;
          16'h164f : blkif.rom_rdata <= 32'h00000000;
          16'h1650 : blkif.rom_rdata <= 32'h00000000;
          16'h1651 : blkif.rom_rdata <= 32'h00000000;
          16'h1652 : blkif.rom_rdata <= 32'h00000000;
          16'h1653 : blkif.rom_rdata <= 32'h00000000;
          16'h1654 : blkif.rom_rdata <= 32'h00000000;
          16'h1655 : blkif.rom_rdata <= 32'h00000000;
          16'h1656 : blkif.rom_rdata <= 32'h00000000;
          16'h1657 : blkif.rom_rdata <= 32'h00000000;
          16'h1658 : blkif.rom_rdata <= 32'h00000000;
          16'h1659 : blkif.rom_rdata <= 32'h00000000;
          16'h165a : blkif.rom_rdata <= 32'h00000000;
          16'h165b : blkif.rom_rdata <= 32'h00000000;
          16'h165c : blkif.rom_rdata <= 32'h00000000;
          16'h165d : blkif.rom_rdata <= 32'h00000000;
          16'h165e : blkif.rom_rdata <= 32'h00000000;
          16'h165f : blkif.rom_rdata <= 32'h00000000;
          16'h1660 : blkif.rom_rdata <= 32'h00000000;
          16'h1661 : blkif.rom_rdata <= 32'h00000000;
          16'h1662 : blkif.rom_rdata <= 32'h00000000;
          16'h1663 : blkif.rom_rdata <= 32'h00000000;
          16'h1664 : blkif.rom_rdata <= 32'h00000000;
          16'h1665 : blkif.rom_rdata <= 32'h00000000;
          16'h1666 : blkif.rom_rdata <= 32'h00000000;
          16'h1667 : blkif.rom_rdata <= 32'h00000000;
          16'h1668 : blkif.rom_rdata <= 32'h00000000;
          16'h1669 : blkif.rom_rdata <= 32'h00000000;
          16'h166a : blkif.rom_rdata <= 32'h00000000;
          16'h166b : blkif.rom_rdata <= 32'h00000000;
          16'h166c : blkif.rom_rdata <= 32'h00000000;
          16'h166d : blkif.rom_rdata <= 32'h00000000;
          16'h166e : blkif.rom_rdata <= 32'h00000000;
          16'h166f : blkif.rom_rdata <= 32'h00000000;
          16'h1670 : blkif.rom_rdata <= 32'h00000000;
          16'h1671 : blkif.rom_rdata <= 32'h00000000;
          16'h1672 : blkif.rom_rdata <= 32'h00000000;
          16'h1673 : blkif.rom_rdata <= 32'h00000000;
          16'h1674 : blkif.rom_rdata <= 32'h00000000;
          16'h1675 : blkif.rom_rdata <= 32'h00000000;
          16'h1676 : blkif.rom_rdata <= 32'h00000000;
          16'h1677 : blkif.rom_rdata <= 32'h00000000;
          16'h1678 : blkif.rom_rdata <= 32'h00000000;
          16'h1679 : blkif.rom_rdata <= 32'h00000000;
          16'h167a : blkif.rom_rdata <= 32'h00000000;
          16'h167b : blkif.rom_rdata <= 32'h00000000;
          16'h167c : blkif.rom_rdata <= 32'h00000000;
          16'h167d : blkif.rom_rdata <= 32'h00000000;
          16'h167e : blkif.rom_rdata <= 32'h00000000;
          16'h167f : blkif.rom_rdata <= 32'h00000000;
          16'h1680 : blkif.rom_rdata <= 32'h00000000;
          16'h1681 : blkif.rom_rdata <= 32'h00000000;
          16'h1682 : blkif.rom_rdata <= 32'h00000000;
          16'h1683 : blkif.rom_rdata <= 32'h00000000;
          16'h1684 : blkif.rom_rdata <= 32'h00000000;
          16'h1685 : blkif.rom_rdata <= 32'h00000000;
          16'h1686 : blkif.rom_rdata <= 32'h00000000;
          16'h1687 : blkif.rom_rdata <= 32'h00000000;
          16'h1688 : blkif.rom_rdata <= 32'h00000000;
          16'h1689 : blkif.rom_rdata <= 32'h00000000;
          16'h168a : blkif.rom_rdata <= 32'h00000000;
          16'h168b : blkif.rom_rdata <= 32'h00000000;
          16'h168c : blkif.rom_rdata <= 32'h00000000;
          16'h168d : blkif.rom_rdata <= 32'h00000000;
          16'h168e : blkif.rom_rdata <= 32'h00000000;
          16'h168f : blkif.rom_rdata <= 32'h00000000;
          16'h1690 : blkif.rom_rdata <= 32'h00000000;
          16'h1691 : blkif.rom_rdata <= 32'h00000000;
          16'h1692 : blkif.rom_rdata <= 32'h00000000;
          16'h1693 : blkif.rom_rdata <= 32'h00000000;
          16'h1694 : blkif.rom_rdata <= 32'h00000000;
          16'h1695 : blkif.rom_rdata <= 32'h00000000;
          16'h1696 : blkif.rom_rdata <= 32'h00000000;
          16'h1697 : blkif.rom_rdata <= 32'h00000000;
          16'h1698 : blkif.rom_rdata <= 32'h00000000;
          16'h1699 : blkif.rom_rdata <= 32'h00000000;
          16'h169a : blkif.rom_rdata <= 32'h00000000;
          16'h169b : blkif.rom_rdata <= 32'h00000000;
          16'h169c : blkif.rom_rdata <= 32'h00000000;
          16'h169d : blkif.rom_rdata <= 32'h00000000;
          16'h169e : blkif.rom_rdata <= 32'h00000000;
          16'h169f : blkif.rom_rdata <= 32'h00000000;
          16'h16a0 : blkif.rom_rdata <= 32'h00000000;
          16'h16a1 : blkif.rom_rdata <= 32'h00000000;
          16'h16a2 : blkif.rom_rdata <= 32'h00000000;
          16'h16a3 : blkif.rom_rdata <= 32'h00000000;
          16'h16a4 : blkif.rom_rdata <= 32'h00000000;
          16'h16a5 : blkif.rom_rdata <= 32'h00000000;
          16'h16a6 : blkif.rom_rdata <= 32'h00000000;
          16'h16a7 : blkif.rom_rdata <= 32'h00000000;
          16'h16a8 : blkif.rom_rdata <= 32'h00000000;
          16'h16a9 : blkif.rom_rdata <= 32'h00000000;
          16'h16aa : blkif.rom_rdata <= 32'h00000000;
          16'h16ab : blkif.rom_rdata <= 32'h00000000;
          16'h16ac : blkif.rom_rdata <= 32'h00000000;
          16'h16ad : blkif.rom_rdata <= 32'h00000000;
          16'h16ae : blkif.rom_rdata <= 32'h00000000;
          16'h16af : blkif.rom_rdata <= 32'h00000000;
          16'h16b0 : blkif.rom_rdata <= 32'h00000000;
          16'h16b1 : blkif.rom_rdata <= 32'h00000000;
          16'h16b2 : blkif.rom_rdata <= 32'h00000000;
          16'h16b3 : blkif.rom_rdata <= 32'h00000000;
          16'h16b4 : blkif.rom_rdata <= 32'h00000000;
          16'h16b5 : blkif.rom_rdata <= 32'h00000000;
          16'h16b6 : blkif.rom_rdata <= 32'h00000000;
          16'h16b7 : blkif.rom_rdata <= 32'h00000000;
          16'h16b8 : blkif.rom_rdata <= 32'h00000000;
          16'h16b9 : blkif.rom_rdata <= 32'h00000000;
          16'h16ba : blkif.rom_rdata <= 32'h00000000;
          16'h16bb : blkif.rom_rdata <= 32'h00000000;
          16'h16bc : blkif.rom_rdata <= 32'h00000000;
          16'h16bd : blkif.rom_rdata <= 32'h00000000;
          16'h16be : blkif.rom_rdata <= 32'h00000000;
          16'h16bf : blkif.rom_rdata <= 32'h00000000;
          16'h16c0 : blkif.rom_rdata <= 32'h00000000;
          16'h16c1 : blkif.rom_rdata <= 32'h00000000;
          16'h16c2 : blkif.rom_rdata <= 32'h00000000;
          16'h16c3 : blkif.rom_rdata <= 32'h00000000;
          16'h16c4 : blkif.rom_rdata <= 32'h00000000;
          16'h16c5 : blkif.rom_rdata <= 32'h00000000;
          16'h16c6 : blkif.rom_rdata <= 32'h00000000;
          16'h16c7 : blkif.rom_rdata <= 32'h00000000;
          16'h16c8 : blkif.rom_rdata <= 32'h00000000;
          16'h16c9 : blkif.rom_rdata <= 32'h00000000;
          16'h16ca : blkif.rom_rdata <= 32'h00000000;
          16'h16cb : blkif.rom_rdata <= 32'h00000000;
          16'h16cc : blkif.rom_rdata <= 32'h00000000;
          16'h16cd : blkif.rom_rdata <= 32'h00000000;
          16'h16ce : blkif.rom_rdata <= 32'h00000000;
          16'h16cf : blkif.rom_rdata <= 32'h00000000;
          16'h16d0 : blkif.rom_rdata <= 32'h00000000;
          16'h16d1 : blkif.rom_rdata <= 32'h00000000;
          16'h16d2 : blkif.rom_rdata <= 32'h00000000;
          16'h16d3 : blkif.rom_rdata <= 32'h00000000;
          16'h16d4 : blkif.rom_rdata <= 32'h00000000;
          16'h16d5 : blkif.rom_rdata <= 32'h00000000;
          16'h16d6 : blkif.rom_rdata <= 32'h00000000;
          16'h16d7 : blkif.rom_rdata <= 32'h00000000;
          16'h16d8 : blkif.rom_rdata <= 32'h00000000;
          16'h16d9 : blkif.rom_rdata <= 32'h00000000;
          16'h16da : blkif.rom_rdata <= 32'h00000000;
          16'h16db : blkif.rom_rdata <= 32'h00000000;
          16'h16dc : blkif.rom_rdata <= 32'h00000000;
          16'h16dd : blkif.rom_rdata <= 32'h00000000;
          16'h16de : blkif.rom_rdata <= 32'h00000000;
          16'h16df : blkif.rom_rdata <= 32'h00000000;
          16'h16e0 : blkif.rom_rdata <= 32'h00000000;
          16'h16e1 : blkif.rom_rdata <= 32'h00000000;
          16'h16e2 : blkif.rom_rdata <= 32'h00000000;
          16'h16e3 : blkif.rom_rdata <= 32'h00000000;
          16'h16e4 : blkif.rom_rdata <= 32'h00000000;
          16'h16e5 : blkif.rom_rdata <= 32'h00000000;
          16'h16e6 : blkif.rom_rdata <= 32'h00000000;
          16'h16e7 : blkif.rom_rdata <= 32'h00000000;
          16'h16e8 : blkif.rom_rdata <= 32'h00000000;
          16'h16e9 : blkif.rom_rdata <= 32'h00000000;
          16'h16ea : blkif.rom_rdata <= 32'h00000000;
          16'h16eb : blkif.rom_rdata <= 32'h00000000;
          16'h16ec : blkif.rom_rdata <= 32'h00000000;
          16'h16ed : blkif.rom_rdata <= 32'h00000000;
          16'h16ee : blkif.rom_rdata <= 32'h00000000;
          16'h16ef : blkif.rom_rdata <= 32'h00000000;
          16'h16f0 : blkif.rom_rdata <= 32'h00000000;
          16'h16f1 : blkif.rom_rdata <= 32'h00000000;
          16'h16f2 : blkif.rom_rdata <= 32'h00000000;
          16'h16f3 : blkif.rom_rdata <= 32'h00000000;
          16'h16f4 : blkif.rom_rdata <= 32'h00000000;
          16'h16f5 : blkif.rom_rdata <= 32'h00000000;
          16'h16f6 : blkif.rom_rdata <= 32'h00000000;
          16'h16f7 : blkif.rom_rdata <= 32'h00000000;
          16'h16f8 : blkif.rom_rdata <= 32'h00000000;
          16'h16f9 : blkif.rom_rdata <= 32'h00000000;
          16'h16fa : blkif.rom_rdata <= 32'h00000000;
          16'h16fb : blkif.rom_rdata <= 32'h00000000;
          16'h16fc : blkif.rom_rdata <= 32'h00000000;
          16'h16fd : blkif.rom_rdata <= 32'h00000000;
          16'h16fe : blkif.rom_rdata <= 32'h00000000;
          16'h16ff : blkif.rom_rdata <= 32'h00000000;
          16'h1700 : blkif.rom_rdata <= 32'h00000000;
          16'h1701 : blkif.rom_rdata <= 32'h00000000;
          16'h1702 : blkif.rom_rdata <= 32'h00000000;
          16'h1703 : blkif.rom_rdata <= 32'h00000000;
          16'h1704 : blkif.rom_rdata <= 32'h00000000;
          16'h1705 : blkif.rom_rdata <= 32'h00000000;
          16'h1706 : blkif.rom_rdata <= 32'h00000000;
          16'h1707 : blkif.rom_rdata <= 32'h00000000;
          16'h1708 : blkif.rom_rdata <= 32'h00000000;
          16'h1709 : blkif.rom_rdata <= 32'h00000000;
          16'h170a : blkif.rom_rdata <= 32'h00000000;
          16'h170b : blkif.rom_rdata <= 32'h00000000;
          16'h170c : blkif.rom_rdata <= 32'h00000000;
          16'h170d : blkif.rom_rdata <= 32'h00000000;
          16'h170e : blkif.rom_rdata <= 32'h00000000;
          16'h170f : blkif.rom_rdata <= 32'h00000000;
          16'h1710 : blkif.rom_rdata <= 32'h00000000;
          16'h1711 : blkif.rom_rdata <= 32'h00000000;
          16'h1712 : blkif.rom_rdata <= 32'h00000000;
          16'h1713 : blkif.rom_rdata <= 32'h00000000;
          16'h1714 : blkif.rom_rdata <= 32'h00000000;
          16'h1715 : blkif.rom_rdata <= 32'h00000000;
          16'h1716 : blkif.rom_rdata <= 32'h00000000;
          16'h1717 : blkif.rom_rdata <= 32'h00000000;
          16'h1718 : blkif.rom_rdata <= 32'h00000000;
          16'h1719 : blkif.rom_rdata <= 32'h00000000;
          16'h171a : blkif.rom_rdata <= 32'h00000000;
          16'h171b : blkif.rom_rdata <= 32'h00000000;
          16'h171c : blkif.rom_rdata <= 32'h00000000;
          16'h171d : blkif.rom_rdata <= 32'h00000000;
          16'h171e : blkif.rom_rdata <= 32'h00000000;
          16'h171f : blkif.rom_rdata <= 32'h00000000;
          16'h1720 : blkif.rom_rdata <= 32'h00000000;
          16'h1721 : blkif.rom_rdata <= 32'h00000000;
          16'h1722 : blkif.rom_rdata <= 32'h00000000;
          16'h1723 : blkif.rom_rdata <= 32'h00000000;
          16'h1724 : blkif.rom_rdata <= 32'h00000000;
          16'h1725 : blkif.rom_rdata <= 32'h00000000;
          16'h1726 : blkif.rom_rdata <= 32'h00000000;
          16'h1727 : blkif.rom_rdata <= 32'h00000000;
          16'h1728 : blkif.rom_rdata <= 32'h00000000;
          16'h1729 : blkif.rom_rdata <= 32'h00000000;
          16'h172a : blkif.rom_rdata <= 32'h00000000;
          16'h172b : blkif.rom_rdata <= 32'h00000000;
          16'h172c : blkif.rom_rdata <= 32'h00000000;
          16'h172d : blkif.rom_rdata <= 32'h00000000;
          16'h172e : blkif.rom_rdata <= 32'h00000000;
          16'h172f : blkif.rom_rdata <= 32'h00000000;
          16'h1730 : blkif.rom_rdata <= 32'h00000000;
          16'h1731 : blkif.rom_rdata <= 32'h00000000;
          16'h1732 : blkif.rom_rdata <= 32'h00000000;
          16'h1733 : blkif.rom_rdata <= 32'h00000000;
          16'h1734 : blkif.rom_rdata <= 32'h00000000;
          16'h1735 : blkif.rom_rdata <= 32'h00000000;
          16'h1736 : blkif.rom_rdata <= 32'h00000000;
          16'h1737 : blkif.rom_rdata <= 32'h00000000;
          16'h1738 : blkif.rom_rdata <= 32'h00000000;
          16'h1739 : blkif.rom_rdata <= 32'h00000000;
          16'h173a : blkif.rom_rdata <= 32'h00000000;
          16'h173b : blkif.rom_rdata <= 32'h00000000;
          16'h173c : blkif.rom_rdata <= 32'h00000000;
          16'h173d : blkif.rom_rdata <= 32'h00000000;
          16'h173e : blkif.rom_rdata <= 32'h00000000;
          16'h173f : blkif.rom_rdata <= 32'h00000000;
          16'h1740 : blkif.rom_rdata <= 32'h00000000;
          16'h1741 : blkif.rom_rdata <= 32'h00000000;
          16'h1742 : blkif.rom_rdata <= 32'h00000000;
          16'h1743 : blkif.rom_rdata <= 32'h00000000;
          16'h1744 : blkif.rom_rdata <= 32'h00000000;
          16'h1745 : blkif.rom_rdata <= 32'h00000000;
          16'h1746 : blkif.rom_rdata <= 32'h00000000;
          16'h1747 : blkif.rom_rdata <= 32'h00000000;
          16'h1748 : blkif.rom_rdata <= 32'h00000000;
          16'h1749 : blkif.rom_rdata <= 32'h00000000;
          16'h174a : blkif.rom_rdata <= 32'h00000000;
          16'h174b : blkif.rom_rdata <= 32'h00000000;
          16'h174c : blkif.rom_rdata <= 32'h00000000;
          16'h174d : blkif.rom_rdata <= 32'h00000000;
          16'h174e : blkif.rom_rdata <= 32'h00000000;
          16'h174f : blkif.rom_rdata <= 32'h00000000;
          16'h1750 : blkif.rom_rdata <= 32'h00000000;
          16'h1751 : blkif.rom_rdata <= 32'h00000000;
          16'h1752 : blkif.rom_rdata <= 32'h00000000;
          16'h1753 : blkif.rom_rdata <= 32'h00000000;
          16'h1754 : blkif.rom_rdata <= 32'h00000000;
          16'h1755 : blkif.rom_rdata <= 32'h00000000;
          16'h1756 : blkif.rom_rdata <= 32'h00000000;
          16'h1757 : blkif.rom_rdata <= 32'h00000000;
          16'h1758 : blkif.rom_rdata <= 32'h00000000;
          16'h1759 : blkif.rom_rdata <= 32'h00000000;
          16'h175a : blkif.rom_rdata <= 32'h00000000;
          16'h175b : blkif.rom_rdata <= 32'h00000000;
          16'h175c : blkif.rom_rdata <= 32'h00000000;
          16'h175d : blkif.rom_rdata <= 32'h00000000;
          16'h175e : blkif.rom_rdata <= 32'h00000000;
          16'h175f : blkif.rom_rdata <= 32'h00000000;
          16'h1760 : blkif.rom_rdata <= 32'h00000000;
          16'h1761 : blkif.rom_rdata <= 32'h00000000;
          16'h1762 : blkif.rom_rdata <= 32'h00000000;
          16'h1763 : blkif.rom_rdata <= 32'h00000000;
          16'h1764 : blkif.rom_rdata <= 32'h00000000;
          16'h1765 : blkif.rom_rdata <= 32'h00000000;
          16'h1766 : blkif.rom_rdata <= 32'h00000000;
          16'h1767 : blkif.rom_rdata <= 32'h00000000;
          16'h1768 : blkif.rom_rdata <= 32'h00000000;
          16'h1769 : blkif.rom_rdata <= 32'h00000000;
          16'h176a : blkif.rom_rdata <= 32'h00000000;
          16'h176b : blkif.rom_rdata <= 32'h00000000;
          16'h176c : blkif.rom_rdata <= 32'h00000000;
          16'h176d : blkif.rom_rdata <= 32'h00000000;
          16'h176e : blkif.rom_rdata <= 32'h00000000;
          16'h176f : blkif.rom_rdata <= 32'h00000000;
          16'h1770 : blkif.rom_rdata <= 32'h00000000;
          16'h1771 : blkif.rom_rdata <= 32'h00000000;
          16'h1772 : blkif.rom_rdata <= 32'h00000000;
          16'h1773 : blkif.rom_rdata <= 32'h00000000;
          16'h1774 : blkif.rom_rdata <= 32'h00000000;
          16'h1775 : blkif.rom_rdata <= 32'h00000000;
          16'h1776 : blkif.rom_rdata <= 32'h00000000;
          16'h1777 : blkif.rom_rdata <= 32'h00000000;
          16'h1778 : blkif.rom_rdata <= 32'h00000000;
          16'h1779 : blkif.rom_rdata <= 32'h00000000;
          16'h177a : blkif.rom_rdata <= 32'h00000000;
          16'h177b : blkif.rom_rdata <= 32'h00000000;
          16'h177c : blkif.rom_rdata <= 32'h00000000;
          16'h177d : blkif.rom_rdata <= 32'h00000000;
          16'h177e : blkif.rom_rdata <= 32'h00000000;
          16'h177f : blkif.rom_rdata <= 32'h00000000;
          16'h1780 : blkif.rom_rdata <= 32'h00000000;
          16'h1781 : blkif.rom_rdata <= 32'h00000000;
          16'h1782 : blkif.rom_rdata <= 32'h00000000;
          16'h1783 : blkif.rom_rdata <= 32'h00000000;
          16'h1784 : blkif.rom_rdata <= 32'h00000000;
          16'h1785 : blkif.rom_rdata <= 32'h00000000;
          16'h1786 : blkif.rom_rdata <= 32'h00000000;
          16'h1787 : blkif.rom_rdata <= 32'h00000000;
          16'h1788 : blkif.rom_rdata <= 32'h00000000;
          16'h1789 : blkif.rom_rdata <= 32'h00000000;
          16'h178a : blkif.rom_rdata <= 32'h00000000;
          16'h178b : blkif.rom_rdata <= 32'h00000000;
          16'h178c : blkif.rom_rdata <= 32'h00000000;
          16'h178d : blkif.rom_rdata <= 32'h00000000;
          16'h178e : blkif.rom_rdata <= 32'h00000000;
          16'h178f : blkif.rom_rdata <= 32'h00000000;
          16'h1790 : blkif.rom_rdata <= 32'h00000000;
          16'h1791 : blkif.rom_rdata <= 32'h00000000;
          16'h1792 : blkif.rom_rdata <= 32'h00000000;
          16'h1793 : blkif.rom_rdata <= 32'h00000000;
          16'h1794 : blkif.rom_rdata <= 32'h00000000;
          16'h1795 : blkif.rom_rdata <= 32'h00000000;
          16'h1796 : blkif.rom_rdata <= 32'h00000000;
          16'h1797 : blkif.rom_rdata <= 32'h00000000;
          16'h1798 : blkif.rom_rdata <= 32'h00000000;
          16'h1799 : blkif.rom_rdata <= 32'h00000000;
          16'h179a : blkif.rom_rdata <= 32'h00000000;
          16'h179b : blkif.rom_rdata <= 32'h00000000;
          16'h179c : blkif.rom_rdata <= 32'h00000000;
          16'h179d : blkif.rom_rdata <= 32'h00000000;
          16'h179e : blkif.rom_rdata <= 32'h00000000;
          16'h179f : blkif.rom_rdata <= 32'h00000000;
          16'h17a0 : blkif.rom_rdata <= 32'h00000000;
          16'h17a1 : blkif.rom_rdata <= 32'h00000000;
          16'h17a2 : blkif.rom_rdata <= 32'h00000000;
          16'h17a3 : blkif.rom_rdata <= 32'h00000000;
          16'h17a4 : blkif.rom_rdata <= 32'h00000000;
          16'h17a5 : blkif.rom_rdata <= 32'h00000000;
          16'h17a6 : blkif.rom_rdata <= 32'h00000000;
          16'h17a7 : blkif.rom_rdata <= 32'h00000000;
          16'h17a8 : blkif.rom_rdata <= 32'h00000000;
          16'h17a9 : blkif.rom_rdata <= 32'h00000000;
          16'h17aa : blkif.rom_rdata <= 32'h00000000;
          16'h17ab : blkif.rom_rdata <= 32'h00000000;
          16'h17ac : blkif.rom_rdata <= 32'h00000000;
          16'h17ad : blkif.rom_rdata <= 32'h00000000;
          16'h17ae : blkif.rom_rdata <= 32'h00000000;
          16'h17af : blkif.rom_rdata <= 32'h00000000;
          16'h17b0 : blkif.rom_rdata <= 32'h00000000;
          16'h17b1 : blkif.rom_rdata <= 32'h00000000;
          16'h17b2 : blkif.rom_rdata <= 32'h00000000;
          16'h17b3 : blkif.rom_rdata <= 32'h00000000;
          16'h17b4 : blkif.rom_rdata <= 32'h00000000;
          16'h17b5 : blkif.rom_rdata <= 32'h00000000;
          16'h17b6 : blkif.rom_rdata <= 32'h00000000;
          16'h17b7 : blkif.rom_rdata <= 32'h00000000;
          16'h17b8 : blkif.rom_rdata <= 32'h00000000;
          16'h17b9 : blkif.rom_rdata <= 32'h00000000;
          16'h17ba : blkif.rom_rdata <= 32'h00000000;
          16'h17bb : blkif.rom_rdata <= 32'h00000000;
          16'h17bc : blkif.rom_rdata <= 32'h00000000;
          16'h17bd : blkif.rom_rdata <= 32'h00000000;
          16'h17be : blkif.rom_rdata <= 32'h00000000;
          16'h17bf : blkif.rom_rdata <= 32'h00000000;
          16'h17c0 : blkif.rom_rdata <= 32'h00000000;
          16'h17c1 : blkif.rom_rdata <= 32'h00000000;
          16'h17c2 : blkif.rom_rdata <= 32'h00000000;
          16'h17c3 : blkif.rom_rdata <= 32'h00000000;
          16'h17c4 : blkif.rom_rdata <= 32'h00000000;
          16'h17c5 : blkif.rom_rdata <= 32'h00000000;
          16'h17c6 : blkif.rom_rdata <= 32'h00000000;
          16'h17c7 : blkif.rom_rdata <= 32'h00000000;
          16'h17c8 : blkif.rom_rdata <= 32'h00000000;
          16'h17c9 : blkif.rom_rdata <= 32'h00000000;
          16'h17ca : blkif.rom_rdata <= 32'h00000000;
          16'h17cb : blkif.rom_rdata <= 32'h00000000;
          16'h17cc : blkif.rom_rdata <= 32'h00000000;
          16'h17cd : blkif.rom_rdata <= 32'h00000000;
          16'h17ce : blkif.rom_rdata <= 32'h00000000;
          16'h17cf : blkif.rom_rdata <= 32'h00000000;
          16'h17d0 : blkif.rom_rdata <= 32'h00000000;
          16'h17d1 : blkif.rom_rdata <= 32'h00000000;
          16'h17d2 : blkif.rom_rdata <= 32'h00000000;
          16'h17d3 : blkif.rom_rdata <= 32'h00000000;
          16'h17d4 : blkif.rom_rdata <= 32'h00000000;
          16'h17d5 : blkif.rom_rdata <= 32'h00000000;
          16'h17d6 : blkif.rom_rdata <= 32'h00000000;
          16'h17d7 : blkif.rom_rdata <= 32'h00000000;
          16'h17d8 : blkif.rom_rdata <= 32'h00000000;
          16'h17d9 : blkif.rom_rdata <= 32'h00000000;
          16'h17da : blkif.rom_rdata <= 32'h00000000;
          16'h17db : blkif.rom_rdata <= 32'h00000000;
          16'h17dc : blkif.rom_rdata <= 32'h00000000;
          16'h17dd : blkif.rom_rdata <= 32'h00000000;
          16'h17de : blkif.rom_rdata <= 32'h00000000;
          16'h17df : blkif.rom_rdata <= 32'h00000000;
          16'h17e0 : blkif.rom_rdata <= 32'h00000000;
          16'h17e1 : blkif.rom_rdata <= 32'h00000000;
          16'h17e2 : blkif.rom_rdata <= 32'h00000000;
          16'h17e3 : blkif.rom_rdata <= 32'h00000000;
          16'h17e4 : blkif.rom_rdata <= 32'h00000000;
          16'h17e5 : blkif.rom_rdata <= 32'h00000000;
          16'h17e6 : blkif.rom_rdata <= 32'h00000000;
          16'h17e7 : blkif.rom_rdata <= 32'h00000000;
          16'h17e8 : blkif.rom_rdata <= 32'h00000000;
          16'h17e9 : blkif.rom_rdata <= 32'h00000000;
          16'h17ea : blkif.rom_rdata <= 32'h00000000;
          16'h17eb : blkif.rom_rdata <= 32'h00000000;
          16'h17ec : blkif.rom_rdata <= 32'h00000000;
          16'h17ed : blkif.rom_rdata <= 32'h00000000;
          16'h17ee : blkif.rom_rdata <= 32'h00000000;
          16'h17ef : blkif.rom_rdata <= 32'h00000000;
          16'h17f0 : blkif.rom_rdata <= 32'h00000000;
          16'h17f1 : blkif.rom_rdata <= 32'h00000000;
          16'h17f2 : blkif.rom_rdata <= 32'h00000000;
          16'h17f3 : blkif.rom_rdata <= 32'h00000000;
          16'h17f4 : blkif.rom_rdata <= 32'h00000000;
          16'h17f5 : blkif.rom_rdata <= 32'h00000000;
          16'h17f6 : blkif.rom_rdata <= 32'h00000000;
          16'h17f7 : blkif.rom_rdata <= 32'h00000000;
          16'h17f8 : blkif.rom_rdata <= 32'h00000000;
          16'h17f9 : blkif.rom_rdata <= 32'h00000000;
          16'h17fa : blkif.rom_rdata <= 32'h00000000;
          16'h17fb : blkif.rom_rdata <= 32'h00000000;
          16'h17fc : blkif.rom_rdata <= 32'h00000000;
          16'h17fd : blkif.rom_rdata <= 32'h00000000;
          16'h17fe : blkif.rom_rdata <= 32'h00000000;
          16'h17ff : blkif.rom_rdata <= 32'h00000000;
          16'h1800 : blkif.rom_rdata <= 32'ha4500000;
          16'h1801 : blkif.rom_rdata <= 32'h24190000;
          16'h1802 : blkif.rom_rdata <= 32'h18510000;
          16'h1803 : blkif.rom_rdata <= 32'h20190000;
          16'h1804 : blkif.rom_rdata <= 32'h18510000;
          16'h1805 : blkif.rom_rdata <= 32'h21190000;
          16'h1806 : blkif.rom_rdata <= 32'h18510000;
          16'h1807 : blkif.rom_rdata <= 32'h22190000;
          16'h1808 : blkif.rom_rdata <= 32'h18510000;
          16'h1809 : blkif.rom_rdata <= 32'h23190000;
          16'h180a : blkif.rom_rdata <= 32'h18510000;
          16'h180b : blkif.rom_rdata <= 32'h24190000;
          16'h180c : blkif.rom_rdata <= 32'h18510000;
          16'h180d : blkif.rom_rdata <= 32'h25190000;
          16'h180e : blkif.rom_rdata <= 32'h18510000;
          16'h180f : blkif.rom_rdata <= 32'h26190000;
          16'h1810 : blkif.rom_rdata <= 32'h18510000;
          16'h1811 : blkif.rom_rdata <= 32'h27190000;
          16'h1812 : blkif.rom_rdata <= 32'h18510000;
          16'h1813 : blkif.rom_rdata <= 32'h28190000;
          16'h1814 : blkif.rom_rdata <= 32'h18510000;
          16'h1815 : blkif.rom_rdata <= 32'h29190000;
          16'h1816 : blkif.rom_rdata <= 32'h18510000;
          16'h1817 : blkif.rom_rdata <= 32'h2a190000;
          16'h1818 : blkif.rom_rdata <= 32'h18510000;
          16'h1819 : blkif.rom_rdata <= 32'h2b190000;
          16'h181a : blkif.rom_rdata <= 32'h18510000;
          16'h181b : blkif.rom_rdata <= 32'h2c190000;
          16'h181c : blkif.rom_rdata <= 32'h18510000;
          16'h181d : blkif.rom_rdata <= 32'h2d190000;
          16'h181e : blkif.rom_rdata <= 32'h18510000;
          16'h181f : blkif.rom_rdata <= 32'h2e190000;
          16'h1820 : blkif.rom_rdata <= 32'h18510000;
          16'h1821 : blkif.rom_rdata <= 32'h2f190000;
          16'h1822 : blkif.rom_rdata <= 32'h18510000;
          16'h1823 : blkif.rom_rdata <= 32'h30190000;
          16'h1824 : blkif.rom_rdata <= 32'h18510000;
          16'h1825 : blkif.rom_rdata <= 32'h31190000;
          16'h1826 : blkif.rom_rdata <= 32'h18510000;
          16'h1827 : blkif.rom_rdata <= 32'h32190000;
          16'h1828 : blkif.rom_rdata <= 32'h18510000;
          16'h1829 : blkif.rom_rdata <= 32'h33190000;
          16'h182a : blkif.rom_rdata <= 32'h18510000;
          16'h182b : blkif.rom_rdata <= 32'h34190000;
          16'h182c : blkif.rom_rdata <= 32'h18510000;
          16'h182d : blkif.rom_rdata <= 32'h35190000;
          16'h182e : blkif.rom_rdata <= 32'h18510000;
          16'h182f : blkif.rom_rdata <= 32'h36190000;
          16'h1830 : blkif.rom_rdata <= 32'h18510000;
          16'h1831 : blkif.rom_rdata <= 32'h37190000;
          16'h1832 : blkif.rom_rdata <= 32'h18510000;
          16'h1833 : blkif.rom_rdata <= 32'h38190000;
          16'h1834 : blkif.rom_rdata <= 32'h18510000;
          16'h1835 : blkif.rom_rdata <= 32'h39190000;
          16'h1836 : blkif.rom_rdata <= 32'h18510000;
          16'h1837 : blkif.rom_rdata <= 32'h3a190000;
          16'h1838 : blkif.rom_rdata <= 32'h18510000;
          16'h1839 : blkif.rom_rdata <= 32'h3b190000;
          16'h183a : blkif.rom_rdata <= 32'h18510000;
          16'h183b : blkif.rom_rdata <= 32'h3c190000;
          16'h183c : blkif.rom_rdata <= 32'h18510000;
          16'h183d : blkif.rom_rdata <= 32'h3d190000;
          16'h183e : blkif.rom_rdata <= 32'h18510000;
          16'h183f : blkif.rom_rdata <= 32'h3e190000;
          16'h1840 : blkif.rom_rdata <= 32'h18510000;
          16'h1841 : blkif.rom_rdata <= 32'h3f190000;
          16'h1842 : blkif.rom_rdata <= 32'h9c520000;
          16'h1843 : blkif.rom_rdata <= 32'h22190000;
          16'h1844 : blkif.rom_rdata <= 32'hb0520000;
          16'h1845 : blkif.rom_rdata <= 32'h22190000;
          16'h1846 : blkif.rom_rdata <= 32'hc0520000;
          16'h1847 : blkif.rom_rdata <= 32'h02190000;
          16'h1848 : blkif.rom_rdata <= 32'hd0520000;
          16'h1849 : blkif.rom_rdata <= 32'h02190000;
          16'h184a : blkif.rom_rdata <= 32'hb0530000;
          16'h184b : blkif.rom_rdata <= 32'h22190000;
          16'h184c : blkif.rom_rdata <= 32'hc0530000;
          16'h184d : blkif.rom_rdata <= 32'h22190000;
          16'h184e : blkif.rom_rdata <= 32'hd4530000;
          16'h184f : blkif.rom_rdata <= 32'h02190000;
          16'h1850 : blkif.rom_rdata <= 32'he8530000;
          16'h1851 : blkif.rom_rdata <= 32'h02190000;
          16'h1852 : blkif.rom_rdata <= 32'h08550000;
          16'h1853 : blkif.rom_rdata <= 32'h22190000;
          16'h1854 : blkif.rom_rdata <= 32'h14550000;
          16'h1855 : blkif.rom_rdata <= 32'h22190000;
          16'h1856 : blkif.rom_rdata <= 32'h28550000;
          16'h1857 : blkif.rom_rdata <= 32'h02190000;
          16'h1858 : blkif.rom_rdata <= 32'h34550000;
          16'h1859 : blkif.rom_rdata <= 32'h02190000;
          16'h185a : blkif.rom_rdata <= 32'h48550000;
          16'h185b : blkif.rom_rdata <= 32'h02190000;
          16'h185c : blkif.rom_rdata <= 32'hfc550000;
          16'h185d : blkif.rom_rdata <= 32'h22190000;
          16'h185e : blkif.rom_rdata <= 32'h08560000;
          16'h185f : blkif.rom_rdata <= 32'h22190000;
          16'h1860 : blkif.rom_rdata <= 32'h1c560000;
          16'h1861 : blkif.rom_rdata <= 32'h02190000;
          16'h1862 : blkif.rom_rdata <= 32'h80560000;
          16'h1863 : blkif.rom_rdata <= 32'h22190000;
          16'h1864 : blkif.rom_rdata <= 32'h18570000;
          16'h1865 : blkif.rom_rdata <= 32'h22190000;
          16'h1866 : blkif.rom_rdata <= 32'h30570000;
          16'h1867 : blkif.rom_rdata <= 32'h02190000;
          16'h1868 : blkif.rom_rdata <= 32'h4c570000;
          16'h1869 : blkif.rom_rdata <= 32'h02190000;
          16'h186a : blkif.rom_rdata <= 32'hff00f00f;
          16'h186b : blkif.rom_rdata <= 32'hff00f00f;
          16'h186c : blkif.rom_rdata <= 32'hff0000ff;
          16'h186d : blkif.rom_rdata <= 32'hf00f0ff0;
          16'h186e : blkif.rom_rdata <= 32'hff0000ff;
          16'h186f : blkif.rom_rdata <= 32'hf00f0ff0;
          16'h1870 : blkif.rom_rdata <= 32'hff00ff00;
          16'h1871 : blkif.rom_rdata <= 32'h00ff00ff;
          16'h1872 : blkif.rom_rdata <= 32'hf00ff00f;
          16'h1873 : blkif.rom_rdata <= 32'h0ff00ff0;
          16'h1874 : blkif.rom_rdata <= 32'h00000000;
          16'h1875 : blkif.rom_rdata <= 32'h00000000;
          16'h1876 : blkif.rom_rdata <= 32'h00000000;
          16'h1877 : blkif.rom_rdata <= 32'h00000000;
          16'h1878 : blkif.rom_rdata <= 32'h00000000;
          16'h1879 : blkif.rom_rdata <= 32'h00000000;
          16'h187a : blkif.rom_rdata <= 32'h00000000;
          16'h187b : blkif.rom_rdata <= 32'h00000000;
          16'h187c : blkif.rom_rdata <= 32'h00000000;
          16'h187d : blkif.rom_rdata <= 32'h00000000;
          16'h187e : blkif.rom_rdata <= 32'h00000000;
          16'h187f : blkif.rom_rdata <= 32'h00000000;
          16'h1880 : blkif.rom_rdata <= 32'h00000000;
          16'h1881 : blkif.rom_rdata <= 32'h00000000;
          16'h1882 : blkif.rom_rdata <= 32'h00000000;
          16'h1883 : blkif.rom_rdata <= 32'h00000000;
          16'h1884 : blkif.rom_rdata <= 32'h00000000;
          16'h1885 : blkif.rom_rdata <= 32'h00000000;
          16'h1886 : blkif.rom_rdata <= 32'h00000000;
          16'h1887 : blkif.rom_rdata <= 32'h00000000;
          16'h1888 : blkif.rom_rdata <= 32'h00000000;
          16'h1889 : blkif.rom_rdata <= 32'h00000000;
          16'h188a : blkif.rom_rdata <= 32'h00000000;
          16'h188b : blkif.rom_rdata <= 32'h00000000;
          16'h188c : blkif.rom_rdata <= 32'h00000000;
          16'h188d : blkif.rom_rdata <= 32'h00000000;
          16'h188e : blkif.rom_rdata <= 32'h00000000;
          16'h188f : blkif.rom_rdata <= 32'h00000000;
          16'h1890 : blkif.rom_rdata <= 32'h00000000;
          16'h1891 : blkif.rom_rdata <= 32'h00000000;
          16'h1892 : blkif.rom_rdata <= 32'h00000000;
          16'h1893 : blkif.rom_rdata <= 32'h00000000;
          16'h1894 : blkif.rom_rdata <= 32'h00000000;
          16'h1895 : blkif.rom_rdata <= 32'h00000000;
          16'h1896 : blkif.rom_rdata <= 32'h00000000;
          16'h1897 : blkif.rom_rdata <= 32'h00000000;
          16'h1898 : blkif.rom_rdata <= 32'h00000000;
          16'h1899 : blkif.rom_rdata <= 32'h00000000;
          16'h189a : blkif.rom_rdata <= 32'h00000000;
          16'h189b : blkif.rom_rdata <= 32'h00000000;
          16'h189c : blkif.rom_rdata <= 32'h00000000;
          16'h189d : blkif.rom_rdata <= 32'h00000000;
          16'h189e : blkif.rom_rdata <= 32'h00000000;
          16'h189f : blkif.rom_rdata <= 32'h00000000;
          16'h18a0 : blkif.rom_rdata <= 32'h00000000;
          16'h18a1 : blkif.rom_rdata <= 32'h00000000;
          16'h18a2 : blkif.rom_rdata <= 32'h00000000;
          16'h18a3 : blkif.rom_rdata <= 32'h00000000;
          16'h18a4 : blkif.rom_rdata <= 32'h00000000;
          16'h18a5 : blkif.rom_rdata <= 32'h00000000;
          16'h18a6 : blkif.rom_rdata <= 32'h00000000;
          16'h18a7 : blkif.rom_rdata <= 32'h00000000;
          16'h18a8 : blkif.rom_rdata <= 32'h00000000;
          16'h18a9 : blkif.rom_rdata <= 32'h00000000;
          16'h18aa : blkif.rom_rdata <= 32'h00000000;
          16'h18ab : blkif.rom_rdata <= 32'h00000000;
          16'h18ac : blkif.rom_rdata <= 32'h00000000;
          16'h18ad : blkif.rom_rdata <= 32'h00000000;
          16'h18ae : blkif.rom_rdata <= 32'h00000000;
          16'h18af : blkif.rom_rdata <= 32'h00000000;
          16'h18b0 : blkif.rom_rdata <= 32'h00000000;
          16'h18b1 : blkif.rom_rdata <= 32'h00000000;
          16'h18b2 : blkif.rom_rdata <= 32'h00000000;
          16'h18b3 : blkif.rom_rdata <= 32'h00000000;
          16'h18b4 : blkif.rom_rdata <= 32'h00000000;
          16'h18b5 : blkif.rom_rdata <= 32'h00000000;
          16'h18b6 : blkif.rom_rdata <= 32'h00000000;
          16'h18b7 : blkif.rom_rdata <= 32'h00000000;
          16'h18b8 : blkif.rom_rdata <= 32'h00000000;
          16'h18b9 : blkif.rom_rdata <= 32'h00000000;
          16'h18ba : blkif.rom_rdata <= 32'h00000000;
          16'h18bb : blkif.rom_rdata <= 32'h00000000;
          16'h18bc : blkif.rom_rdata <= 32'h00000000;
          16'h18bd : blkif.rom_rdata <= 32'h00000000;
          16'h18be : blkif.rom_rdata <= 32'h00000000;
          16'h18bf : blkif.rom_rdata <= 32'h00000000;
          16'h18c0 : blkif.rom_rdata <= 32'h00000000;
          16'h18c1 : blkif.rom_rdata <= 32'h00000000;
          16'h18c2 : blkif.rom_rdata <= 32'h00000000;
          16'h18c3 : blkif.rom_rdata <= 32'h00000000;
          16'h18c4 : blkif.rom_rdata <= 32'h00000000;
          16'h18c5 : blkif.rom_rdata <= 32'h00000000;
          16'h18c6 : blkif.rom_rdata <= 32'h00000000;
          16'h18c7 : blkif.rom_rdata <= 32'h00000000;
          16'h18c8 : blkif.rom_rdata <= 32'h00000000;
          16'h18c9 : blkif.rom_rdata <= 32'h00000000;
          16'h18ca : blkif.rom_rdata <= 32'h00000000;
          16'h18cb : blkif.rom_rdata <= 32'h00000000;
          16'h18cc : blkif.rom_rdata <= 32'h00000000;
          16'h18cd : blkif.rom_rdata <= 32'h00000000;
          16'h18ce : blkif.rom_rdata <= 32'h00000000;
          16'h18cf : blkif.rom_rdata <= 32'h00000000;
          16'h18d0 : blkif.rom_rdata <= 32'h00000000;
          16'h18d1 : blkif.rom_rdata <= 32'h00000000;
          16'h18d2 : blkif.rom_rdata <= 32'h00000000;
          16'h18d3 : blkif.rom_rdata <= 32'h00000000;
          16'h18d4 : blkif.rom_rdata <= 32'h00000000;
          16'h18d5 : blkif.rom_rdata <= 32'h00000000;
          16'h18d6 : blkif.rom_rdata <= 32'h00000000;
          16'h18d7 : blkif.rom_rdata <= 32'h00000000;
          16'h18d8 : blkif.rom_rdata <= 32'h00000000;
          16'h18d9 : blkif.rom_rdata <= 32'h00000000;
          16'h18da : blkif.rom_rdata <= 32'h00000000;
          16'h18db : blkif.rom_rdata <= 32'h00000000;
          16'h18dc : blkif.rom_rdata <= 32'h00000000;
          16'h18dd : blkif.rom_rdata <= 32'h00000000;
          16'h18de : blkif.rom_rdata <= 32'h00000000;
          16'h18df : blkif.rom_rdata <= 32'h00000000;
          16'h18e0 : blkif.rom_rdata <= 32'h00000000;
          16'h18e1 : blkif.rom_rdata <= 32'h00000000;
          16'h18e2 : blkif.rom_rdata <= 32'h00000000;
          16'h18e3 : blkif.rom_rdata <= 32'h00000000;
          16'h18e4 : blkif.rom_rdata <= 32'h00000000;
          16'h18e5 : blkif.rom_rdata <= 32'h00000000;
          16'h18e6 : blkif.rom_rdata <= 32'h00000000;
          16'h18e7 : blkif.rom_rdata <= 32'h00000000;
          16'h18e8 : blkif.rom_rdata <= 32'h00000000;
          16'h18e9 : blkif.rom_rdata <= 32'h00000000;
          16'h18ea : blkif.rom_rdata <= 32'h00000000;
          16'h18eb : blkif.rom_rdata <= 32'h00000000;
          16'h18ec : blkif.rom_rdata <= 32'h00000000;
          16'h18ed : blkif.rom_rdata <= 32'h00000000;
          16'h18ee : blkif.rom_rdata <= 32'h00000000;
          16'h18ef : blkif.rom_rdata <= 32'h00000000;
          16'h18f0 : blkif.rom_rdata <= 32'h00000000;
          16'h18f1 : blkif.rom_rdata <= 32'h00000000;
          16'h18f2 : blkif.rom_rdata <= 32'h00000000;
          16'h18f3 : blkif.rom_rdata <= 32'h00000000;
          16'h18f4 : blkif.rom_rdata <= 32'h00000000;
          16'h18f5 : blkif.rom_rdata <= 32'h00000000;
          16'h18f6 : blkif.rom_rdata <= 32'h00000000;
          16'h18f7 : blkif.rom_rdata <= 32'h00000000;
          16'h18f8 : blkif.rom_rdata <= 32'h00000000;
          16'h18f9 : blkif.rom_rdata <= 32'h00000000;
          16'h18fa : blkif.rom_rdata <= 32'h00000000;
          16'h18fb : blkif.rom_rdata <= 32'h00000000;
          16'h18fc : blkif.rom_rdata <= 32'h00000000;
          16'h18fd : blkif.rom_rdata <= 32'h00000000;
          16'h18fe : blkif.rom_rdata <= 32'h00000000;
          16'h18ff : blkif.rom_rdata <= 32'h00000000;
          16'h1900 : blkif.rom_rdata <= 32'h00000000;
          16'h1901 : blkif.rom_rdata <= 32'h00000000;
          16'h1902 : blkif.rom_rdata <= 32'h00000000;
          16'h1903 : blkif.rom_rdata <= 32'h00000000;
          16'h1904 : blkif.rom_rdata <= 32'h00000000;
          16'h1905 : blkif.rom_rdata <= 32'h00000000;
          16'h1906 : blkif.rom_rdata <= 32'h00000000;
          16'h1907 : blkif.rom_rdata <= 32'h00000000;
          16'h1908 : blkif.rom_rdata <= 32'h00000000;
          16'h1909 : blkif.rom_rdata <= 32'h00000000;
          16'h190a : blkif.rom_rdata <= 32'h00000000;
          16'h190b : blkif.rom_rdata <= 32'h00000000;
          16'h190c : blkif.rom_rdata <= 32'h00000000;
          16'h190d : blkif.rom_rdata <= 32'h00000000;
          16'h190e : blkif.rom_rdata <= 32'h00000000;
          16'h190f : blkif.rom_rdata <= 32'h00000000;
          16'h1910 : blkif.rom_rdata <= 32'h00000000;
          16'h1911 : blkif.rom_rdata <= 32'h00000000;
          16'h1912 : blkif.rom_rdata <= 32'h00000000;
          16'h1913 : blkif.rom_rdata <= 32'h00000000;
          16'h1914 : blkif.rom_rdata <= 32'h00000000;
          16'h1915 : blkif.rom_rdata <= 32'h00000000;
          16'h1916 : blkif.rom_rdata <= 32'h00000000;
          16'h1917 : blkif.rom_rdata <= 32'h00000000;
          16'h1918 : blkif.rom_rdata <= 32'h00000000;
          16'h1919 : blkif.rom_rdata <= 32'h00000000;
          16'h191a : blkif.rom_rdata <= 32'h00000000;
          16'h191b : blkif.rom_rdata <= 32'h00000000;
          16'h191c : blkif.rom_rdata <= 32'h00000000;
          16'h191d : blkif.rom_rdata <= 32'h00000000;
          16'h191e : blkif.rom_rdata <= 32'h00000000;
          16'h191f : blkif.rom_rdata <= 32'h00000000;
          16'h1920 : blkif.rom_rdata <= 32'h00000000;
          16'h1921 : blkif.rom_rdata <= 32'h00000000;
          16'h1922 : blkif.rom_rdata <= 32'h00000000;
          16'h1923 : blkif.rom_rdata <= 32'h00000000;
          16'h1924 : blkif.rom_rdata <= 32'h00000000;
          16'h1925 : blkif.rom_rdata <= 32'h00000000;
          16'h1926 : blkif.rom_rdata <= 32'h00000000;
          16'h1927 : blkif.rom_rdata <= 32'h00000000;
          16'h1928 : blkif.rom_rdata <= 32'h00000000;
          16'h1929 : blkif.rom_rdata <= 32'h00000000;
          16'h192a : blkif.rom_rdata <= 32'h00000000;
          16'h192b : blkif.rom_rdata <= 32'h00000000;
          16'h192c : blkif.rom_rdata <= 32'h00000000;
          16'h192d : blkif.rom_rdata <= 32'h00000000;
          16'h192e : blkif.rom_rdata <= 32'h00000000;
          16'h192f : blkif.rom_rdata <= 32'h00000000;
          16'h1930 : blkif.rom_rdata <= 32'h00000000;
          16'h1931 : blkif.rom_rdata <= 32'h00000000;
          16'h1932 : blkif.rom_rdata <= 32'h00000000;
          16'h1933 : blkif.rom_rdata <= 32'h00000000;
          16'h1934 : blkif.rom_rdata <= 32'h00000000;
          16'h1935 : blkif.rom_rdata <= 32'h00000000;
          16'h1936 : blkif.rom_rdata <= 32'h00000000;
          16'h1937 : blkif.rom_rdata <= 32'h00000000;
          16'h1938 : blkif.rom_rdata <= 32'h00000000;
          16'h1939 : blkif.rom_rdata <= 32'h00000000;
          16'h193a : blkif.rom_rdata <= 32'h00000000;
          16'h193b : blkif.rom_rdata <= 32'h00000000;
          16'h193c : blkif.rom_rdata <= 32'h00000000;
          16'h193d : blkif.rom_rdata <= 32'h00000000;
          16'h193e : blkif.rom_rdata <= 32'h00000000;
          16'h193f : blkif.rom_rdata <= 32'h00000000;
          16'h1940 : blkif.rom_rdata <= 32'h00000000;
          16'h1941 : blkif.rom_rdata <= 32'h00000000;
          16'h1942 : blkif.rom_rdata <= 32'h00000000;
          16'h1943 : blkif.rom_rdata <= 32'h00000000;
          16'h1944 : blkif.rom_rdata <= 32'h00000000;
          16'h1945 : blkif.rom_rdata <= 32'h00000000;
          16'h1946 : blkif.rom_rdata <= 32'h00000000;
          16'h1947 : blkif.rom_rdata <= 32'h00000000;
          16'h1948 : blkif.rom_rdata <= 32'h00000000;
          16'h1949 : blkif.rom_rdata <= 32'h00000000;
          16'h194a : blkif.rom_rdata <= 32'h00000000;
          16'h194b : blkif.rom_rdata <= 32'h00000000;
          16'h194c : blkif.rom_rdata <= 32'h00000000;
          16'h194d : blkif.rom_rdata <= 32'h00000000;
          16'h194e : blkif.rom_rdata <= 32'h00000000;
          16'h194f : blkif.rom_rdata <= 32'h00000000;
          16'h1950 : blkif.rom_rdata <= 32'h00000000;
          16'h1951 : blkif.rom_rdata <= 32'h00000000;
          16'h1952 : blkif.rom_rdata <= 32'h00000000;
          16'h1953 : blkif.rom_rdata <= 32'h00000000;
          16'h1954 : blkif.rom_rdata <= 32'h00000000;
          16'h1955 : blkif.rom_rdata <= 32'h00000000;
          16'h1956 : blkif.rom_rdata <= 32'h00000000;
          16'h1957 : blkif.rom_rdata <= 32'h00000000;
          16'h1958 : blkif.rom_rdata <= 32'h00000000;
          16'h1959 : blkif.rom_rdata <= 32'h00000000;
          16'h195a : blkif.rom_rdata <= 32'h00000000;
          16'h195b : blkif.rom_rdata <= 32'h00000000;
          16'h195c : blkif.rom_rdata <= 32'h00000000;
          16'h195d : blkif.rom_rdata <= 32'h00000000;
          16'h195e : blkif.rom_rdata <= 32'h00000000;
          16'h195f : blkif.rom_rdata <= 32'h00000000;
          16'h1960 : blkif.rom_rdata <= 32'h00000000;
          16'h1961 : blkif.rom_rdata <= 32'h00000000;
          16'h1962 : blkif.rom_rdata <= 32'h00000000;
          16'h1963 : blkif.rom_rdata <= 32'h00000000;
          16'h1964 : blkif.rom_rdata <= 32'h00000000;
          16'h1965 : blkif.rom_rdata <= 32'h00000000;
          16'h1966 : blkif.rom_rdata <= 32'h00000000;
          16'h1967 : blkif.rom_rdata <= 32'h00000000;
          16'h1968 : blkif.rom_rdata <= 32'h00000000;
          16'h1969 : blkif.rom_rdata <= 32'h00000000;
          16'h196a : blkif.rom_rdata <= 32'h00000000;
          16'h196b : blkif.rom_rdata <= 32'h00000000;
          16'h196c : blkif.rom_rdata <= 32'h00000000;
          16'h196d : blkif.rom_rdata <= 32'h00000000;
          16'h196e : blkif.rom_rdata <= 32'h00000000;
          16'h196f : blkif.rom_rdata <= 32'h00000000;
          16'h1970 : blkif.rom_rdata <= 32'h00000000;
          16'h1971 : blkif.rom_rdata <= 32'h00000000;
          16'h1972 : blkif.rom_rdata <= 32'h00000000;
          16'h1973 : blkif.rom_rdata <= 32'h00000000;
          16'h1974 : blkif.rom_rdata <= 32'h00000000;
          16'h1975 : blkif.rom_rdata <= 32'h00000000;
          16'h1976 : blkif.rom_rdata <= 32'h00000000;
          16'h1977 : blkif.rom_rdata <= 32'h00000000;
          16'h1978 : blkif.rom_rdata <= 32'h00000000;
          16'h1979 : blkif.rom_rdata <= 32'h00000000;
          16'h197a : blkif.rom_rdata <= 32'h00000000;
          16'h197b : blkif.rom_rdata <= 32'h00000000;
          16'h197c : blkif.rom_rdata <= 32'h00000000;
          16'h197d : blkif.rom_rdata <= 32'h00000000;
          16'h197e : blkif.rom_rdata <= 32'h00000000;
          16'h197f : blkif.rom_rdata <= 32'h00000000;
          16'h1980 : blkif.rom_rdata <= 32'h00000000;
          16'h1981 : blkif.rom_rdata <= 32'h00000000;
          16'h1982 : blkif.rom_rdata <= 32'h00000000;
          16'h1983 : blkif.rom_rdata <= 32'h00000000;
          16'h1984 : blkif.rom_rdata <= 32'h00000000;
          16'h1985 : blkif.rom_rdata <= 32'h00000000;
          16'h1986 : blkif.rom_rdata <= 32'h00000000;
          16'h1987 : blkif.rom_rdata <= 32'h00000000;
          16'h1988 : blkif.rom_rdata <= 32'h00000000;
          16'h1989 : blkif.rom_rdata <= 32'h00000000;
          16'h198a : blkif.rom_rdata <= 32'h00000000;
          16'h198b : blkif.rom_rdata <= 32'h00000000;
          16'h198c : blkif.rom_rdata <= 32'h00000000;
          16'h198d : blkif.rom_rdata <= 32'h00000000;
          16'h198e : blkif.rom_rdata <= 32'h00000000;
          16'h198f : blkif.rom_rdata <= 32'h00000000;
          16'h1990 : blkif.rom_rdata <= 32'h00000000;
          16'h1991 : blkif.rom_rdata <= 32'h00000000;
          16'h1992 : blkif.rom_rdata <= 32'h00000000;
          16'h1993 : blkif.rom_rdata <= 32'h00000000;
          16'h1994 : blkif.rom_rdata <= 32'h00000000;
          16'h1995 : blkif.rom_rdata <= 32'h00000000;
          16'h1996 : blkif.rom_rdata <= 32'h00000000;
          16'h1997 : blkif.rom_rdata <= 32'h00000000;
          16'h1998 : blkif.rom_rdata <= 32'h00000000;
          16'h1999 : blkif.rom_rdata <= 32'h00000000;
          16'h199a : blkif.rom_rdata <= 32'h00000000;
          16'h199b : blkif.rom_rdata <= 32'h00000000;
          16'h199c : blkif.rom_rdata <= 32'h00000000;
          16'h199d : blkif.rom_rdata <= 32'h00000000;
          16'h199e : blkif.rom_rdata <= 32'h00000000;
          16'h199f : blkif.rom_rdata <= 32'h00000000;
          16'h19a0 : blkif.rom_rdata <= 32'h00000000;
          16'h19a1 : blkif.rom_rdata <= 32'h00000000;
          16'h19a2 : blkif.rom_rdata <= 32'h00000000;
          16'h19a3 : blkif.rom_rdata <= 32'h00000000;
          16'h19a4 : blkif.rom_rdata <= 32'h00000000;
          16'h19a5 : blkif.rom_rdata <= 32'h00000000;
          16'h19a6 : blkif.rom_rdata <= 32'h00000000;
          16'h19a7 : blkif.rom_rdata <= 32'h00000000;
          16'h19a8 : blkif.rom_rdata <= 32'h00000000;
          16'h19a9 : blkif.rom_rdata <= 32'h00000000;
          16'h19aa : blkif.rom_rdata <= 32'h00000000;
          16'h19ab : blkif.rom_rdata <= 32'h00000000;
          16'h19ac : blkif.rom_rdata <= 32'h00000000;
          16'h19ad : blkif.rom_rdata <= 32'h00000000;
          16'h19ae : blkif.rom_rdata <= 32'h00000000;
          16'h19af : blkif.rom_rdata <= 32'h00000000;
          16'h19b0 : blkif.rom_rdata <= 32'h00000000;
          16'h19b1 : blkif.rom_rdata <= 32'h00000000;
          16'h19b2 : blkif.rom_rdata <= 32'h00000000;
          16'h19b3 : blkif.rom_rdata <= 32'h00000000;
          16'h19b4 : blkif.rom_rdata <= 32'h00000000;
          16'h19b5 : blkif.rom_rdata <= 32'h00000000;
          16'h19b6 : blkif.rom_rdata <= 32'h00000000;
          16'h19b7 : blkif.rom_rdata <= 32'h00000000;
          16'h19b8 : blkif.rom_rdata <= 32'h00000000;
          16'h19b9 : blkif.rom_rdata <= 32'h00000000;
          16'h19ba : blkif.rom_rdata <= 32'h00000000;
          16'h19bb : blkif.rom_rdata <= 32'h00000000;
          16'h19bc : blkif.rom_rdata <= 32'h00000000;
          16'h19bd : blkif.rom_rdata <= 32'h00000000;
          16'h19be : blkif.rom_rdata <= 32'h00000000;
          16'h19bf : blkif.rom_rdata <= 32'h00000000;
          16'h19c0 : blkif.rom_rdata <= 32'h00000000;
          16'h19c1 : blkif.rom_rdata <= 32'h00000000;
          16'h19c2 : blkif.rom_rdata <= 32'h00000000;
          16'h19c3 : blkif.rom_rdata <= 32'h00000000;
          16'h19c4 : blkif.rom_rdata <= 32'h00000000;
          16'h19c5 : blkif.rom_rdata <= 32'h00000000;
          16'h19c6 : blkif.rom_rdata <= 32'h00000000;
          16'h19c7 : blkif.rom_rdata <= 32'h00000000;
          16'h19c8 : blkif.rom_rdata <= 32'h00000000;
          16'h19c9 : blkif.rom_rdata <= 32'h00000000;
          16'h19ca : blkif.rom_rdata <= 32'h00000000;
          16'h19cb : blkif.rom_rdata <= 32'h00000000;
          16'h19cc : blkif.rom_rdata <= 32'h00000000;
          16'h19cd : blkif.rom_rdata <= 32'h00000000;
          16'h19ce : blkif.rom_rdata <= 32'h00000000;
          16'h19cf : blkif.rom_rdata <= 32'h00000000;
          16'h19d0 : blkif.rom_rdata <= 32'h00000000;
          16'h19d1 : blkif.rom_rdata <= 32'h00000000;
          16'h19d2 : blkif.rom_rdata <= 32'h00000000;
          16'h19d3 : blkif.rom_rdata <= 32'h00000000;
          16'h19d4 : blkif.rom_rdata <= 32'h00000000;
          16'h19d5 : blkif.rom_rdata <= 32'h00000000;
          16'h19d6 : blkif.rom_rdata <= 32'h00000000;
          16'h19d7 : blkif.rom_rdata <= 32'h00000000;
          16'h19d8 : blkif.rom_rdata <= 32'h00000000;
          16'h19d9 : blkif.rom_rdata <= 32'h00000000;
          16'h19da : blkif.rom_rdata <= 32'h00000000;
          16'h19db : blkif.rom_rdata <= 32'h00000000;
          16'h19dc : blkif.rom_rdata <= 32'h00000000;
          16'h19dd : blkif.rom_rdata <= 32'h00000000;
          16'h19de : blkif.rom_rdata <= 32'h00000000;
          16'h19df : blkif.rom_rdata <= 32'h00000000;
          16'h19e0 : blkif.rom_rdata <= 32'h00000000;
          16'h19e1 : blkif.rom_rdata <= 32'h00000000;
          16'h19e2 : blkif.rom_rdata <= 32'h00000000;
          16'h19e3 : blkif.rom_rdata <= 32'h00000000;
          16'h19e4 : blkif.rom_rdata <= 32'h00000000;
          16'h19e5 : blkif.rom_rdata <= 32'h00000000;
          16'h19e6 : blkif.rom_rdata <= 32'h00000000;
          16'h19e7 : blkif.rom_rdata <= 32'h00000000;
          16'h19e8 : blkif.rom_rdata <= 32'h00000000;
          16'h19e9 : blkif.rom_rdata <= 32'h00000000;
          16'h19ea : blkif.rom_rdata <= 32'h00000000;
          16'h19eb : blkif.rom_rdata <= 32'h00000000;
          16'h19ec : blkif.rom_rdata <= 32'h00000000;
          16'h19ed : blkif.rom_rdata <= 32'h00000000;
          16'h19ee : blkif.rom_rdata <= 32'h00000000;
          16'h19ef : blkif.rom_rdata <= 32'h00000000;
          16'h19f0 : blkif.rom_rdata <= 32'h00000000;
          16'h19f1 : blkif.rom_rdata <= 32'h00000000;
          16'h19f2 : blkif.rom_rdata <= 32'h00000000;
          16'h19f3 : blkif.rom_rdata <= 32'h00000000;
          16'h19f4 : blkif.rom_rdata <= 32'h00000000;
          16'h19f5 : blkif.rom_rdata <= 32'h00000000;
          16'h19f6 : blkif.rom_rdata <= 32'h00000000;
          16'h19f7 : blkif.rom_rdata <= 32'h00000000;
          16'h19f8 : blkif.rom_rdata <= 32'h00000000;
          16'h19f9 : blkif.rom_rdata <= 32'h00000000;
          16'h19fa : blkif.rom_rdata <= 32'h00000000;
          16'h19fb : blkif.rom_rdata <= 32'h00000000;
          16'h19fc : blkif.rom_rdata <= 32'h00000000;
          16'h19fd : blkif.rom_rdata <= 32'h00000000;
          16'h19fe : blkif.rom_rdata <= 32'h00000000;
          16'h19ff : blkif.rom_rdata <= 32'h00000000;
          16'h1a00 : blkif.rom_rdata <= 32'h00000000;
          16'h1a01 : blkif.rom_rdata <= 32'h00000000;
          16'h1a02 : blkif.rom_rdata <= 32'h00000000;
          16'h1a03 : blkif.rom_rdata <= 32'h00000000;
          16'h1a04 : blkif.rom_rdata <= 32'h00000000;
          16'h1a05 : blkif.rom_rdata <= 32'h00000000;
          16'h1a06 : blkif.rom_rdata <= 32'h00000000;
          16'h1a07 : blkif.rom_rdata <= 32'h00000000;
          16'h1a08 : blkif.rom_rdata <= 32'h00000000;
          16'h1a09 : blkif.rom_rdata <= 32'h00000000;
          16'h1a0a : blkif.rom_rdata <= 32'h00000000;
          16'h1a0b : blkif.rom_rdata <= 32'h00000000;
          16'h1a0c : blkif.rom_rdata <= 32'h00000000;
          16'h1a0d : blkif.rom_rdata <= 32'h00000000;
          16'h1a0e : blkif.rom_rdata <= 32'h00000000;
          16'h1a0f : blkif.rom_rdata <= 32'h00000000;
          16'h1a10 : blkif.rom_rdata <= 32'h00000000;
          16'h1a11 : blkif.rom_rdata <= 32'h00000000;
          16'h1a12 : blkif.rom_rdata <= 32'h00000000;
          16'h1a13 : blkif.rom_rdata <= 32'h00000000;
          16'h1a14 : blkif.rom_rdata <= 32'h00000000;
          16'h1a15 : blkif.rom_rdata <= 32'h00000000;
          16'h1a16 : blkif.rom_rdata <= 32'h00000000;
          16'h1a17 : blkif.rom_rdata <= 32'h00000000;
          16'h1a18 : blkif.rom_rdata <= 32'h00000000;
          16'h1a19 : blkif.rom_rdata <= 32'h00000000;
          16'h1a1a : blkif.rom_rdata <= 32'h00000000;
          16'h1a1b : blkif.rom_rdata <= 32'h00000000;
          16'h1a1c : blkif.rom_rdata <= 32'h00000000;
          16'h1a1d : blkif.rom_rdata <= 32'h00000000;
          16'h1a1e : blkif.rom_rdata <= 32'h00000000;
          16'h1a1f : blkif.rom_rdata <= 32'h00000000;
          16'h1a20 : blkif.rom_rdata <= 32'h00000000;
          16'h1a21 : blkif.rom_rdata <= 32'h00000000;
          16'h1a22 : blkif.rom_rdata <= 32'h00000000;
          16'h1a23 : blkif.rom_rdata <= 32'h00000000;
          16'h1a24 : blkif.rom_rdata <= 32'h00000000;
          16'h1a25 : blkif.rom_rdata <= 32'h00000000;
          16'h1a26 : blkif.rom_rdata <= 32'h00000000;
          16'h1a27 : blkif.rom_rdata <= 32'h00000000;
          16'h1a28 : blkif.rom_rdata <= 32'h00000000;
          16'h1a29 : blkif.rom_rdata <= 32'h00000000;
          16'h1a2a : blkif.rom_rdata <= 32'h00000000;
          16'h1a2b : blkif.rom_rdata <= 32'h00000000;
          16'h1a2c : blkif.rom_rdata <= 32'h00000000;
          16'h1a2d : blkif.rom_rdata <= 32'h00000000;
          16'h1a2e : blkif.rom_rdata <= 32'h00000000;
          16'h1a2f : blkif.rom_rdata <= 32'h00000000;
          16'h1a30 : blkif.rom_rdata <= 32'h00000000;
          16'h1a31 : blkif.rom_rdata <= 32'h00000000;
          16'h1a32 : blkif.rom_rdata <= 32'h00000000;
          16'h1a33 : blkif.rom_rdata <= 32'h00000000;
          16'h1a34 : blkif.rom_rdata <= 32'h00000000;
          16'h1a35 : blkif.rom_rdata <= 32'h00000000;
          16'h1a36 : blkif.rom_rdata <= 32'h00000000;
          16'h1a37 : blkif.rom_rdata <= 32'h00000000;
          16'h1a38 : blkif.rom_rdata <= 32'h00000000;
          16'h1a39 : blkif.rom_rdata <= 32'h00000000;
          16'h1a3a : blkif.rom_rdata <= 32'h00000000;
          16'h1a3b : blkif.rom_rdata <= 32'h00000000;
          16'h1a3c : blkif.rom_rdata <= 32'h00000000;
          16'h1a3d : blkif.rom_rdata <= 32'h00000000;
          16'h1a3e : blkif.rom_rdata <= 32'h00000000;
          16'h1a3f : blkif.rom_rdata <= 32'h00000000;
          16'h1a40 : blkif.rom_rdata <= 32'h00000000;
          16'h1a41 : blkif.rom_rdata <= 32'h00000000;
          16'h1a42 : blkif.rom_rdata <= 32'h00000000;
          16'h1a43 : blkif.rom_rdata <= 32'h00000000;
          16'h1a44 : blkif.rom_rdata <= 32'h00000000;
          16'h1a45 : blkif.rom_rdata <= 32'h00000000;
          16'h1a46 : blkif.rom_rdata <= 32'h00000000;
          16'h1a47 : blkif.rom_rdata <= 32'h00000000;
          16'h1a48 : blkif.rom_rdata <= 32'h00000000;
          16'h1a49 : blkif.rom_rdata <= 32'h00000000;
          16'h1a4a : blkif.rom_rdata <= 32'h00000000;
          16'h1a4b : blkif.rom_rdata <= 32'h00000000;
          16'h1a4c : blkif.rom_rdata <= 32'h00000000;
          16'h1a4d : blkif.rom_rdata <= 32'h00000000;
          16'h1a4e : blkif.rom_rdata <= 32'h00000000;
          16'h1a4f : blkif.rom_rdata <= 32'h00000000;
          16'h1a50 : blkif.rom_rdata <= 32'h00000000;
          16'h1a51 : blkif.rom_rdata <= 32'h00000000;
          16'h1a52 : blkif.rom_rdata <= 32'h00000000;
          16'h1a53 : blkif.rom_rdata <= 32'h00000000;
          16'h1a54 : blkif.rom_rdata <= 32'h00000000;
          16'h1a55 : blkif.rom_rdata <= 32'h00000000;
          16'h1a56 : blkif.rom_rdata <= 32'h00000000;
          16'h1a57 : blkif.rom_rdata <= 32'h00000000;
          16'h1a58 : blkif.rom_rdata <= 32'h00000000;
          16'h1a59 : blkif.rom_rdata <= 32'h00000000;
          16'h1a5a : blkif.rom_rdata <= 32'h00000000;
          16'h1a5b : blkif.rom_rdata <= 32'h00000000;
          16'h1a5c : blkif.rom_rdata <= 32'h00000000;
          16'h1a5d : blkif.rom_rdata <= 32'h00000000;
          16'h1a5e : blkif.rom_rdata <= 32'h00000000;
          16'h1a5f : blkif.rom_rdata <= 32'h00000000;
          16'h1a60 : blkif.rom_rdata <= 32'h00000000;
          16'h1a61 : blkif.rom_rdata <= 32'h00000000;
          16'h1a62 : blkif.rom_rdata <= 32'h00000000;
          16'h1a63 : blkif.rom_rdata <= 32'h00000000;
          16'h1a64 : blkif.rom_rdata <= 32'h00000000;
          16'h1a65 : blkif.rom_rdata <= 32'h00000000;
          16'h1a66 : blkif.rom_rdata <= 32'h00000000;
          16'h1a67 : blkif.rom_rdata <= 32'h00000000;
          16'h1a68 : blkif.rom_rdata <= 32'h00000000;
          16'h1a69 : blkif.rom_rdata <= 32'h00000000;
          16'h1a6a : blkif.rom_rdata <= 32'h00000000;
          16'h1a6b : blkif.rom_rdata <= 32'h00000000;
          16'h1a6c : blkif.rom_rdata <= 32'h00000000;
          16'h1a6d : blkif.rom_rdata <= 32'h00000000;
          16'h1a6e : blkif.rom_rdata <= 32'h00000000;
          16'h1a6f : blkif.rom_rdata <= 32'h00000000;
          16'h1a70 : blkif.rom_rdata <= 32'h00000000;
          16'h1a71 : blkif.rom_rdata <= 32'h00000000;
          16'h1a72 : blkif.rom_rdata <= 32'h00000000;
          16'h1a73 : blkif.rom_rdata <= 32'h00000000;
          16'h1a74 : blkif.rom_rdata <= 32'h00000000;
          16'h1a75 : blkif.rom_rdata <= 32'h00000000;
          16'h1a76 : blkif.rom_rdata <= 32'h00000000;
          16'h1a77 : blkif.rom_rdata <= 32'h00000000;
          16'h1a78 : blkif.rom_rdata <= 32'h00000000;
          16'h1a79 : blkif.rom_rdata <= 32'h00000000;
          16'h1a7a : blkif.rom_rdata <= 32'h00000000;
          16'h1a7b : blkif.rom_rdata <= 32'h00000000;
          16'h1a7c : blkif.rom_rdata <= 32'h00000000;
          16'h1a7d : blkif.rom_rdata <= 32'h00000000;
          16'h1a7e : blkif.rom_rdata <= 32'h00000000;
          16'h1a7f : blkif.rom_rdata <= 32'h00000000;
          16'h1a80 : blkif.rom_rdata <= 32'h00000000;
          16'h1a81 : blkif.rom_rdata <= 32'h00000000;
          16'h1a82 : blkif.rom_rdata <= 32'h00000000;
          16'h1a83 : blkif.rom_rdata <= 32'h00000000;
          16'h1a84 : blkif.rom_rdata <= 32'h00000000;
          16'h1a85 : blkif.rom_rdata <= 32'h00000000;
          16'h1a86 : blkif.rom_rdata <= 32'h00000000;
          16'h1a87 : blkif.rom_rdata <= 32'h00000000;
          16'h1a88 : blkif.rom_rdata <= 32'h00000000;
          16'h1a89 : blkif.rom_rdata <= 32'h00000000;
          16'h1a8a : blkif.rom_rdata <= 32'h00000000;
          16'h1a8b : blkif.rom_rdata <= 32'h00000000;
          16'h1a8c : blkif.rom_rdata <= 32'h00000000;
          16'h1a8d : blkif.rom_rdata <= 32'h00000000;
          16'h1a8e : blkif.rom_rdata <= 32'h00000000;
          16'h1a8f : blkif.rom_rdata <= 32'h00000000;
          16'h1a90 : blkif.rom_rdata <= 32'h00000000;
          16'h1a91 : blkif.rom_rdata <= 32'h00000000;
          16'h1a92 : blkif.rom_rdata <= 32'h00000000;
          16'h1a93 : blkif.rom_rdata <= 32'h00000000;
          16'h1a94 : blkif.rom_rdata <= 32'h00000000;
          16'h1a95 : blkif.rom_rdata <= 32'h00000000;
          16'h1a96 : blkif.rom_rdata <= 32'h00000000;
          16'h1a97 : blkif.rom_rdata <= 32'h00000000;
          16'h1a98 : blkif.rom_rdata <= 32'h00000000;
          16'h1a99 : blkif.rom_rdata <= 32'h00000000;
          16'h1a9a : blkif.rom_rdata <= 32'h00000000;
          16'h1a9b : blkif.rom_rdata <= 32'h00000000;
          16'h1a9c : blkif.rom_rdata <= 32'h00000000;
          16'h1a9d : blkif.rom_rdata <= 32'h00000000;
          16'h1a9e : blkif.rom_rdata <= 32'h00000000;
          16'h1a9f : blkif.rom_rdata <= 32'h00000000;
          16'h1aa0 : blkif.rom_rdata <= 32'h00000000;
          16'h1aa1 : blkif.rom_rdata <= 32'h00000000;
          16'h1aa2 : blkif.rom_rdata <= 32'h00000000;
          16'h1aa3 : blkif.rom_rdata <= 32'h00000000;
          16'h1aa4 : blkif.rom_rdata <= 32'h00000000;
          16'h1aa5 : blkif.rom_rdata <= 32'h00000000;
          16'h1aa6 : blkif.rom_rdata <= 32'h00000000;
          16'h1aa7 : blkif.rom_rdata <= 32'h00000000;
          16'h1aa8 : blkif.rom_rdata <= 32'h00000000;
          16'h1aa9 : blkif.rom_rdata <= 32'h00000000;
          16'h1aaa : blkif.rom_rdata <= 32'h00000000;
          16'h1aab : blkif.rom_rdata <= 32'h00000000;
          16'h1aac : blkif.rom_rdata <= 32'h00000000;
          16'h1aad : blkif.rom_rdata <= 32'h00000000;
          16'h1aae : blkif.rom_rdata <= 32'h00000000;
          16'h1aaf : blkif.rom_rdata <= 32'h00000000;
          16'h1ab0 : blkif.rom_rdata <= 32'h00000000;
          16'h1ab1 : blkif.rom_rdata <= 32'h00000000;
          16'h1ab2 : blkif.rom_rdata <= 32'h00000000;
          16'h1ab3 : blkif.rom_rdata <= 32'h00000000;
          16'h1ab4 : blkif.rom_rdata <= 32'h00000000;
          16'h1ab5 : blkif.rom_rdata <= 32'h00000000;
          16'h1ab6 : blkif.rom_rdata <= 32'h00000000;
          16'h1ab7 : blkif.rom_rdata <= 32'h00000000;
          16'h1ab8 : blkif.rom_rdata <= 32'h00000000;
          16'h1ab9 : blkif.rom_rdata <= 32'h00000000;
          16'h1aba : blkif.rom_rdata <= 32'h00000000;
          16'h1abb : blkif.rom_rdata <= 32'h00000000;
          16'h1abc : blkif.rom_rdata <= 32'h00000000;
          16'h1abd : blkif.rom_rdata <= 32'h00000000;
          16'h1abe : blkif.rom_rdata <= 32'h00000000;
          16'h1abf : blkif.rom_rdata <= 32'h00000000;
          16'h1ac0 : blkif.rom_rdata <= 32'h00000000;
          16'h1ac1 : blkif.rom_rdata <= 32'h00000000;
          16'h1ac2 : blkif.rom_rdata <= 32'h00000000;
          16'h1ac3 : blkif.rom_rdata <= 32'h00000000;
          16'h1ac4 : blkif.rom_rdata <= 32'h00000000;
          16'h1ac5 : blkif.rom_rdata <= 32'h00000000;
          16'h1ac6 : blkif.rom_rdata <= 32'h00000000;
          16'h1ac7 : blkif.rom_rdata <= 32'h00000000;
          16'h1ac8 : blkif.rom_rdata <= 32'h00000000;
          16'h1ac9 : blkif.rom_rdata <= 32'h00000000;
          16'h1aca : blkif.rom_rdata <= 32'h00000000;
          16'h1acb : blkif.rom_rdata <= 32'h00000000;
          16'h1acc : blkif.rom_rdata <= 32'h00000000;
          16'h1acd : blkif.rom_rdata <= 32'h00000000;
          16'h1ace : blkif.rom_rdata <= 32'h00000000;
          16'h1acf : blkif.rom_rdata <= 32'h00000000;
          16'h1ad0 : blkif.rom_rdata <= 32'h00000000;
          16'h1ad1 : blkif.rom_rdata <= 32'h00000000;
          16'h1ad2 : blkif.rom_rdata <= 32'h00000000;
          16'h1ad3 : blkif.rom_rdata <= 32'h00000000;
          16'h1ad4 : blkif.rom_rdata <= 32'h00000000;
          16'h1ad5 : blkif.rom_rdata <= 32'h00000000;
          16'h1ad6 : blkif.rom_rdata <= 32'h00000000;
          16'h1ad7 : blkif.rom_rdata <= 32'h00000000;
          16'h1ad8 : blkif.rom_rdata <= 32'h00000000;
          16'h1ad9 : blkif.rom_rdata <= 32'h00000000;
          16'h1ada : blkif.rom_rdata <= 32'h00000000;
          16'h1adb : blkif.rom_rdata <= 32'h00000000;
          16'h1adc : blkif.rom_rdata <= 32'h00000000;
          16'h1add : blkif.rom_rdata <= 32'h00000000;
          16'h1ade : blkif.rom_rdata <= 32'h00000000;
          16'h1adf : blkif.rom_rdata <= 32'h00000000;
          16'h1ae0 : blkif.rom_rdata <= 32'h00000000;
          16'h1ae1 : blkif.rom_rdata <= 32'h00000000;
          16'h1ae2 : blkif.rom_rdata <= 32'h00000000;
          16'h1ae3 : blkif.rom_rdata <= 32'h00000000;
          16'h1ae4 : blkif.rom_rdata <= 32'h00000000;
          16'h1ae5 : blkif.rom_rdata <= 32'h00000000;
          16'h1ae6 : blkif.rom_rdata <= 32'h00000000;
          16'h1ae7 : blkif.rom_rdata <= 32'h00000000;
          16'h1ae8 : blkif.rom_rdata <= 32'h00000000;
          16'h1ae9 : blkif.rom_rdata <= 32'h00000000;
          16'h1aea : blkif.rom_rdata <= 32'h00000000;
          16'h1aeb : blkif.rom_rdata <= 32'h00000000;
          16'h1aec : blkif.rom_rdata <= 32'h00000000;
          16'h1aed : blkif.rom_rdata <= 32'h00000000;
          16'h1aee : blkif.rom_rdata <= 32'h00000000;
          16'h1aef : blkif.rom_rdata <= 32'h00000000;
          16'h1af0 : blkif.rom_rdata <= 32'h00000000;
          16'h1af1 : blkif.rom_rdata <= 32'h00000000;
          16'h1af2 : blkif.rom_rdata <= 32'h00000000;
          16'h1af3 : blkif.rom_rdata <= 32'h00000000;
          16'h1af4 : blkif.rom_rdata <= 32'h00000000;
          16'h1af5 : blkif.rom_rdata <= 32'h00000000;
          16'h1af6 : blkif.rom_rdata <= 32'h00000000;
          16'h1af7 : blkif.rom_rdata <= 32'h00000000;
          16'h1af8 : blkif.rom_rdata <= 32'h00000000;
          16'h1af9 : blkif.rom_rdata <= 32'h00000000;
          16'h1afa : blkif.rom_rdata <= 32'h00000000;
          16'h1afb : blkif.rom_rdata <= 32'h00000000;
          16'h1afc : blkif.rom_rdata <= 32'h00000000;
          16'h1afd : blkif.rom_rdata <= 32'h00000000;
          16'h1afe : blkif.rom_rdata <= 32'h00000000;
          16'h1aff : blkif.rom_rdata <= 32'h00000000;
          16'h1b00 : blkif.rom_rdata <= 32'h00000000;
          16'h1b01 : blkif.rom_rdata <= 32'h00000000;
          16'h1b02 : blkif.rom_rdata <= 32'h00000000;
          16'h1b03 : blkif.rom_rdata <= 32'h00000000;
          16'h1b04 : blkif.rom_rdata <= 32'h00000000;
          16'h1b05 : blkif.rom_rdata <= 32'h00000000;
          16'h1b06 : blkif.rom_rdata <= 32'h00000000;
          16'h1b07 : blkif.rom_rdata <= 32'h00000000;
          16'h1b08 : blkif.rom_rdata <= 32'h00000000;
          16'h1b09 : blkif.rom_rdata <= 32'h00000000;
          16'h1b0a : blkif.rom_rdata <= 32'h00000000;
          16'h1b0b : blkif.rom_rdata <= 32'h00000000;
          16'h1b0c : blkif.rom_rdata <= 32'h00000000;
          16'h1b0d : blkif.rom_rdata <= 32'h00000000;
          16'h1b0e : blkif.rom_rdata <= 32'h00000000;
          16'h1b0f : blkif.rom_rdata <= 32'h00000000;
          16'h1b10 : blkif.rom_rdata <= 32'h00000000;
          16'h1b11 : blkif.rom_rdata <= 32'h00000000;
          16'h1b12 : blkif.rom_rdata <= 32'h00000000;
          16'h1b13 : blkif.rom_rdata <= 32'h00000000;
          16'h1b14 : blkif.rom_rdata <= 32'h00000000;
          16'h1b15 : blkif.rom_rdata <= 32'h00000000;
          16'h1b16 : blkif.rom_rdata <= 32'h00000000;
          16'h1b17 : blkif.rom_rdata <= 32'h00000000;
          16'h1b18 : blkif.rom_rdata <= 32'h00000000;
          16'h1b19 : blkif.rom_rdata <= 32'h00000000;
          16'h1b1a : blkif.rom_rdata <= 32'h00000000;
          16'h1b1b : blkif.rom_rdata <= 32'h00000000;
          16'h1b1c : blkif.rom_rdata <= 32'h00000000;
          16'h1b1d : blkif.rom_rdata <= 32'h00000000;
          16'h1b1e : blkif.rom_rdata <= 32'h00000000;
          16'h1b1f : blkif.rom_rdata <= 32'h00000000;
          16'h1b20 : blkif.rom_rdata <= 32'h00000000;
          16'h1b21 : blkif.rom_rdata <= 32'h00000000;
          16'h1b22 : blkif.rom_rdata <= 32'h00000000;
          16'h1b23 : blkif.rom_rdata <= 32'h00000000;
          16'h1b24 : blkif.rom_rdata <= 32'h00000000;
          16'h1b25 : blkif.rom_rdata <= 32'h00000000;
          16'h1b26 : blkif.rom_rdata <= 32'h00000000;
          16'h1b27 : blkif.rom_rdata <= 32'h00000000;
          16'h1b28 : blkif.rom_rdata <= 32'h00000000;
          16'h1b29 : blkif.rom_rdata <= 32'h00000000;
          16'h1b2a : blkif.rom_rdata <= 32'h00000000;
          16'h1b2b : blkif.rom_rdata <= 32'h00000000;
          16'h1b2c : blkif.rom_rdata <= 32'h00000000;
          16'h1b2d : blkif.rom_rdata <= 32'h00000000;
          16'h1b2e : blkif.rom_rdata <= 32'h00000000;
          16'h1b2f : blkif.rom_rdata <= 32'h00000000;
          16'h1b30 : blkif.rom_rdata <= 32'h00000000;
          16'h1b31 : blkif.rom_rdata <= 32'h00000000;
          16'h1b32 : blkif.rom_rdata <= 32'h00000000;
          16'h1b33 : blkif.rom_rdata <= 32'h00000000;
          16'h1b34 : blkif.rom_rdata <= 32'h00000000;
          16'h1b35 : blkif.rom_rdata <= 32'h00000000;
          16'h1b36 : blkif.rom_rdata <= 32'h00000000;
          16'h1b37 : blkif.rom_rdata <= 32'h00000000;
          16'h1b38 : blkif.rom_rdata <= 32'h00000000;
          16'h1b39 : blkif.rom_rdata <= 32'h00000000;
          16'h1b3a : blkif.rom_rdata <= 32'h00000000;
          16'h1b3b : blkif.rom_rdata <= 32'h00000000;
          16'h1b3c : blkif.rom_rdata <= 32'h00000000;
          16'h1b3d : blkif.rom_rdata <= 32'h00000000;
          16'h1b3e : blkif.rom_rdata <= 32'h00000000;
          16'h1b3f : blkif.rom_rdata <= 32'h00000000;
          16'h1b40 : blkif.rom_rdata <= 32'h00000000;
          16'h1b41 : blkif.rom_rdata <= 32'h00000000;
          16'h1b42 : blkif.rom_rdata <= 32'h00000000;
          16'h1b43 : blkif.rom_rdata <= 32'h00000000;
          16'h1b44 : blkif.rom_rdata <= 32'h00000000;
          16'h1b45 : blkif.rom_rdata <= 32'h00000000;
          16'h1b46 : blkif.rom_rdata <= 32'h00000000;
          16'h1b47 : blkif.rom_rdata <= 32'h00000000;
          16'h1b48 : blkif.rom_rdata <= 32'h00000000;
          16'h1b49 : blkif.rom_rdata <= 32'h00000000;
          16'h1b4a : blkif.rom_rdata <= 32'h00000000;
          16'h1b4b : blkif.rom_rdata <= 32'h00000000;
          16'h1b4c : blkif.rom_rdata <= 32'h00000000;
          16'h1b4d : blkif.rom_rdata <= 32'h00000000;
          16'h1b4e : blkif.rom_rdata <= 32'h00000000;
          16'h1b4f : blkif.rom_rdata <= 32'h00000000;
          16'h1b50 : blkif.rom_rdata <= 32'h00000000;
          16'h1b51 : blkif.rom_rdata <= 32'h00000000;
          16'h1b52 : blkif.rom_rdata <= 32'h00000000;
          16'h1b53 : blkif.rom_rdata <= 32'h00000000;
          16'h1b54 : blkif.rom_rdata <= 32'h00000000;
          16'h1b55 : blkif.rom_rdata <= 32'h00000000;
          16'h1b56 : blkif.rom_rdata <= 32'h00000000;
          16'h1b57 : blkif.rom_rdata <= 32'h00000000;
          16'h1b58 : blkif.rom_rdata <= 32'h00000000;
          16'h1b59 : blkif.rom_rdata <= 32'h00000000;
          16'h1b5a : blkif.rom_rdata <= 32'h00000000;
          16'h1b5b : blkif.rom_rdata <= 32'h00000000;
          16'h1b5c : blkif.rom_rdata <= 32'h00000000;
          16'h1b5d : blkif.rom_rdata <= 32'h00000000;
          16'h1b5e : blkif.rom_rdata <= 32'h00000000;
          16'h1b5f : blkif.rom_rdata <= 32'h00000000;
          16'h1b60 : blkif.rom_rdata <= 32'h00000000;
          16'h1b61 : blkif.rom_rdata <= 32'h00000000;
          16'h1b62 : blkif.rom_rdata <= 32'h00000000;
          16'h1b63 : blkif.rom_rdata <= 32'h00000000;
          16'h1b64 : blkif.rom_rdata <= 32'h00000000;
          16'h1b65 : blkif.rom_rdata <= 32'h00000000;
          16'h1b66 : blkif.rom_rdata <= 32'h00000000;
          16'h1b67 : blkif.rom_rdata <= 32'h00000000;
          16'h1b68 : blkif.rom_rdata <= 32'h00000000;
          16'h1b69 : blkif.rom_rdata <= 32'h00000000;
          16'h1b6a : blkif.rom_rdata <= 32'h00000000;
          16'h1b6b : blkif.rom_rdata <= 32'h00000000;
          16'h1b6c : blkif.rom_rdata <= 32'h00000000;
          16'h1b6d : blkif.rom_rdata <= 32'h00000000;
          16'h1b6e : blkif.rom_rdata <= 32'h00000000;
          16'h1b6f : blkif.rom_rdata <= 32'h00000000;
          16'h1b70 : blkif.rom_rdata <= 32'h00000000;
          16'h1b71 : blkif.rom_rdata <= 32'h00000000;
          16'h1b72 : blkif.rom_rdata <= 32'h00000000;
          16'h1b73 : blkif.rom_rdata <= 32'h00000000;
          16'h1b74 : blkif.rom_rdata <= 32'h00000000;
          16'h1b75 : blkif.rom_rdata <= 32'h00000000;
          16'h1b76 : blkif.rom_rdata <= 32'h00000000;
          16'h1b77 : blkif.rom_rdata <= 32'h00000000;
          16'h1b78 : blkif.rom_rdata <= 32'h00000000;
          16'h1b79 : blkif.rom_rdata <= 32'h00000000;
          16'h1b7a : blkif.rom_rdata <= 32'h00000000;
          16'h1b7b : blkif.rom_rdata <= 32'h00000000;
          16'h1b7c : blkif.rom_rdata <= 32'h00000000;
          16'h1b7d : blkif.rom_rdata <= 32'h00000000;
          16'h1b7e : blkif.rom_rdata <= 32'h00000000;
          16'h1b7f : blkif.rom_rdata <= 32'h00000000;
          16'h1b80 : blkif.rom_rdata <= 32'h00000000;
          16'h1b81 : blkif.rom_rdata <= 32'h00000000;
          16'h1b82 : blkif.rom_rdata <= 32'h00000000;
          16'h1b83 : blkif.rom_rdata <= 32'h00000000;
          16'h1b84 : blkif.rom_rdata <= 32'h00000000;
          16'h1b85 : blkif.rom_rdata <= 32'h00000000;
          16'h1b86 : blkif.rom_rdata <= 32'h00000000;
          16'h1b87 : blkif.rom_rdata <= 32'h00000000;
          16'h1b88 : blkif.rom_rdata <= 32'h00000000;
          16'h1b89 : blkif.rom_rdata <= 32'h00000000;
          16'h1b8a : blkif.rom_rdata <= 32'h00000000;
          16'h1b8b : blkif.rom_rdata <= 32'h00000000;
          16'h1b8c : blkif.rom_rdata <= 32'h00000000;
          16'h1b8d : blkif.rom_rdata <= 32'h00000000;
          16'h1b8e : blkif.rom_rdata <= 32'h00000000;
          16'h1b8f : blkif.rom_rdata <= 32'h00000000;
          16'h1b90 : blkif.rom_rdata <= 32'h00000000;
          16'h1b91 : blkif.rom_rdata <= 32'h00000000;
          16'h1b92 : blkif.rom_rdata <= 32'h00000000;
          16'h1b93 : blkif.rom_rdata <= 32'h00000000;
          16'h1b94 : blkif.rom_rdata <= 32'h00000000;
          16'h1b95 : blkif.rom_rdata <= 32'h00000000;
          16'h1b96 : blkif.rom_rdata <= 32'h00000000;
          16'h1b97 : blkif.rom_rdata <= 32'h00000000;
          16'h1b98 : blkif.rom_rdata <= 32'h00000000;
          16'h1b99 : blkif.rom_rdata <= 32'h00000000;
          16'h1b9a : blkif.rom_rdata <= 32'h00000000;
          16'h1b9b : blkif.rom_rdata <= 32'h00000000;
          16'h1b9c : blkif.rom_rdata <= 32'h00000000;
          16'h1b9d : blkif.rom_rdata <= 32'h00000000;
          16'h1b9e : blkif.rom_rdata <= 32'h00000000;
          16'h1b9f : blkif.rom_rdata <= 32'h00000000;
          16'h1ba0 : blkif.rom_rdata <= 32'h00000000;
          16'h1ba1 : blkif.rom_rdata <= 32'h00000000;
          16'h1ba2 : blkif.rom_rdata <= 32'h00000000;
          16'h1ba3 : blkif.rom_rdata <= 32'h00000000;
          16'h1ba4 : blkif.rom_rdata <= 32'h00000000;
          16'h1ba5 : blkif.rom_rdata <= 32'h00000000;
          16'h1ba6 : blkif.rom_rdata <= 32'h00000000;
          16'h1ba7 : blkif.rom_rdata <= 32'h00000000;
          16'h1ba8 : blkif.rom_rdata <= 32'h00000000;
          16'h1ba9 : blkif.rom_rdata <= 32'h00000000;
          16'h1baa : blkif.rom_rdata <= 32'h00000000;
          16'h1bab : blkif.rom_rdata <= 32'h00000000;
          16'h1bac : blkif.rom_rdata <= 32'h00000000;
          16'h1bad : blkif.rom_rdata <= 32'h00000000;
          16'h1bae : blkif.rom_rdata <= 32'h00000000;
          16'h1baf : blkif.rom_rdata <= 32'h00000000;
          16'h1bb0 : blkif.rom_rdata <= 32'h00000000;
          16'h1bb1 : blkif.rom_rdata <= 32'h00000000;
          16'h1bb2 : blkif.rom_rdata <= 32'h00000000;
          16'h1bb3 : blkif.rom_rdata <= 32'h00000000;
          16'h1bb4 : blkif.rom_rdata <= 32'h00000000;
          16'h1bb5 : blkif.rom_rdata <= 32'h00000000;
          16'h1bb6 : blkif.rom_rdata <= 32'h00000000;
          16'h1bb7 : blkif.rom_rdata <= 32'h00000000;
          16'h1bb8 : blkif.rom_rdata <= 32'h00000000;
          16'h1bb9 : blkif.rom_rdata <= 32'h00000000;
          16'h1bba : blkif.rom_rdata <= 32'h00000000;
          16'h1bbb : blkif.rom_rdata <= 32'h00000000;
          16'h1bbc : blkif.rom_rdata <= 32'h00000000;
          16'h1bbd : blkif.rom_rdata <= 32'h00000000;
          16'h1bbe : blkif.rom_rdata <= 32'h00000000;
          16'h1bbf : blkif.rom_rdata <= 32'h00000000;
          16'h1bc0 : blkif.rom_rdata <= 32'h00000000;
          16'h1bc1 : blkif.rom_rdata <= 32'h00000000;
          16'h1bc2 : blkif.rom_rdata <= 32'h00000000;
          16'h1bc3 : blkif.rom_rdata <= 32'h00000000;
          16'h1bc4 : blkif.rom_rdata <= 32'h00000000;
          16'h1bc5 : blkif.rom_rdata <= 32'h00000000;
          16'h1bc6 : blkif.rom_rdata <= 32'h00000000;
          16'h1bc7 : blkif.rom_rdata <= 32'h00000000;
          16'h1bc8 : blkif.rom_rdata <= 32'h00000000;
          16'h1bc9 : blkif.rom_rdata <= 32'h00000000;
          16'h1bca : blkif.rom_rdata <= 32'h00000000;
          16'h1bcb : blkif.rom_rdata <= 32'h00000000;
          16'h1bcc : blkif.rom_rdata <= 32'h00000000;
          16'h1bcd : blkif.rom_rdata <= 32'h00000000;
          16'h1bce : blkif.rom_rdata <= 32'h00000000;
          16'h1bcf : blkif.rom_rdata <= 32'h00000000;
          16'h1bd0 : blkif.rom_rdata <= 32'h00000000;
          16'h1bd1 : blkif.rom_rdata <= 32'h00000000;
          16'h1bd2 : blkif.rom_rdata <= 32'h00000000;
          16'h1bd3 : blkif.rom_rdata <= 32'h00000000;
          16'h1bd4 : blkif.rom_rdata <= 32'h00000000;
          16'h1bd5 : blkif.rom_rdata <= 32'h00000000;
          16'h1bd6 : blkif.rom_rdata <= 32'h00000000;
          16'h1bd7 : blkif.rom_rdata <= 32'h00000000;
          16'h1bd8 : blkif.rom_rdata <= 32'h00000000;
          16'h1bd9 : blkif.rom_rdata <= 32'h00000000;
          16'h1bda : blkif.rom_rdata <= 32'h00000000;
          16'h1bdb : blkif.rom_rdata <= 32'h00000000;
          16'h1bdc : blkif.rom_rdata <= 32'h00000000;
          16'h1bdd : blkif.rom_rdata <= 32'h00000000;
          16'h1bde : blkif.rom_rdata <= 32'h00000000;
          16'h1bdf : blkif.rom_rdata <= 32'h00000000;
          16'h1be0 : blkif.rom_rdata <= 32'h00000000;
          16'h1be1 : blkif.rom_rdata <= 32'h00000000;
          16'h1be2 : blkif.rom_rdata <= 32'h00000000;
          16'h1be3 : blkif.rom_rdata <= 32'h00000000;
          16'h1be4 : blkif.rom_rdata <= 32'h00000000;
          16'h1be5 : blkif.rom_rdata <= 32'h00000000;
          16'h1be6 : blkif.rom_rdata <= 32'h00000000;
          16'h1be7 : blkif.rom_rdata <= 32'h00000000;
          16'h1be8 : blkif.rom_rdata <= 32'h00000000;
          16'h1be9 : blkif.rom_rdata <= 32'h00000000;
          16'h1bea : blkif.rom_rdata <= 32'h00000000;
          16'h1beb : blkif.rom_rdata <= 32'h00000000;
          16'h1bec : blkif.rom_rdata <= 32'h00000000;
          16'h1bed : blkif.rom_rdata <= 32'h00000000;
          16'h1bee : blkif.rom_rdata <= 32'h00000000;
          16'h1bef : blkif.rom_rdata <= 32'h00000000;
          16'h1bf0 : blkif.rom_rdata <= 32'h00000000;
          16'h1bf1 : blkif.rom_rdata <= 32'h00000000;
          16'h1bf2 : blkif.rom_rdata <= 32'h00000000;
          16'h1bf3 : blkif.rom_rdata <= 32'h00000000;
          16'h1bf4 : blkif.rom_rdata <= 32'h00000000;
          16'h1bf5 : blkif.rom_rdata <= 32'h00000000;
          16'h1bf6 : blkif.rom_rdata <= 32'h00000000;
          16'h1bf7 : blkif.rom_rdata <= 32'h00000000;
          16'h1bf8 : blkif.rom_rdata <= 32'h00000000;
          16'h1bf9 : blkif.rom_rdata <= 32'h00000000;
          16'h1bfa : blkif.rom_rdata <= 32'h00000000;
          16'h1bfb : blkif.rom_rdata <= 32'h00000000;
          16'h1bfc : blkif.rom_rdata <= 32'h00000000;
          16'h1bfd : blkif.rom_rdata <= 32'h00000000;
          16'h1bfe : blkif.rom_rdata <= 32'h00000000;
          16'h1bff : blkif.rom_rdata <= 32'h00000000;
          16'h1c00 : blkif.rom_rdata <= 32'h00000000;
          16'h1c01 : blkif.rom_rdata <= 32'h00000000;
          16'h1c02 : blkif.rom_rdata <= 32'h00000000;
          16'h1c03 : blkif.rom_rdata <= 32'h00000000;
          16'h1c04 : blkif.rom_rdata <= 32'h00000000;
          16'h1c05 : blkif.rom_rdata <= 32'h00000000;
          16'h1c06 : blkif.rom_rdata <= 32'h00000000;
          16'h1c07 : blkif.rom_rdata <= 32'h00000000;
          16'h1c08 : blkif.rom_rdata <= 32'h00000000;
          16'h1c09 : blkif.rom_rdata <= 32'h00000000;
          16'h1c0a : blkif.rom_rdata <= 32'h00000000;
          16'h1c0b : blkif.rom_rdata <= 32'h00000000;
          16'h1c0c : blkif.rom_rdata <= 32'h00000000;
          16'h1c0d : blkif.rom_rdata <= 32'h00000000;
          16'h1c0e : blkif.rom_rdata <= 32'h00000000;
          16'h1c0f : blkif.rom_rdata <= 32'h00000000;
          16'h1c10 : blkif.rom_rdata <= 32'h00000000;
          16'h1c11 : blkif.rom_rdata <= 32'h00000000;
          16'h1c12 : blkif.rom_rdata <= 32'h00000000;
          16'h1c13 : blkif.rom_rdata <= 32'h00000000;
          16'h1c14 : blkif.rom_rdata <= 32'h00000000;
          16'h1c15 : blkif.rom_rdata <= 32'h00000000;
          16'h1c16 : blkif.rom_rdata <= 32'h00000000;
          16'h1c17 : blkif.rom_rdata <= 32'h00000000;
          16'h1c18 : blkif.rom_rdata <= 32'h00000000;
          16'h1c19 : blkif.rom_rdata <= 32'h00000000;
          16'h1c1a : blkif.rom_rdata <= 32'h00000000;
          16'h1c1b : blkif.rom_rdata <= 32'h00000000;
          16'h1c1c : blkif.rom_rdata <= 32'h00000000;
          16'h1c1d : blkif.rom_rdata <= 32'h00000000;
          16'h1c1e : blkif.rom_rdata <= 32'h00000000;
          16'h1c1f : blkif.rom_rdata <= 32'h00000000;
          16'h1c20 : blkif.rom_rdata <= 32'h00000000;
          16'h1c21 : blkif.rom_rdata <= 32'h00000000;
          16'h1c22 : blkif.rom_rdata <= 32'h00000000;
          16'h1c23 : blkif.rom_rdata <= 32'h00000000;
          16'h1c24 : blkif.rom_rdata <= 32'h00000000;
          16'h1c25 : blkif.rom_rdata <= 32'h00000000;
          16'h1c26 : blkif.rom_rdata <= 32'h00000000;
          16'h1c27 : blkif.rom_rdata <= 32'h00000000;
          16'h1c28 : blkif.rom_rdata <= 32'h00000000;
          16'h1c29 : blkif.rom_rdata <= 32'h00000000;
          16'h1c2a : blkif.rom_rdata <= 32'h00000000;
          16'h1c2b : blkif.rom_rdata <= 32'h00000000;
          16'h1c2c : blkif.rom_rdata <= 32'h00000000;
          16'h1c2d : blkif.rom_rdata <= 32'h00000000;
          16'h1c2e : blkif.rom_rdata <= 32'h00000000;
          16'h1c2f : blkif.rom_rdata <= 32'h00000000;
          16'h1c30 : blkif.rom_rdata <= 32'h00000000;
          16'h1c31 : blkif.rom_rdata <= 32'h00000000;
          16'h1c32 : blkif.rom_rdata <= 32'h00000000;
          16'h1c33 : blkif.rom_rdata <= 32'h00000000;
          16'h1c34 : blkif.rom_rdata <= 32'h00000000;
          16'h1c35 : blkif.rom_rdata <= 32'h00000000;
          16'h1c36 : blkif.rom_rdata <= 32'h00000000;
          16'h1c37 : blkif.rom_rdata <= 32'h00000000;
          16'h1c38 : blkif.rom_rdata <= 32'h00000000;
          16'h1c39 : blkif.rom_rdata <= 32'h00000000;
          16'h1c3a : blkif.rom_rdata <= 32'h00000000;
          16'h1c3b : blkif.rom_rdata <= 32'h00000000;
          16'h1c3c : blkif.rom_rdata <= 32'h00000000;
          16'h1c3d : blkif.rom_rdata <= 32'h00000000;
          16'h1c3e : blkif.rom_rdata <= 32'h00000000;
          16'h1c3f : blkif.rom_rdata <= 32'h00000000;
          16'h1c40 : blkif.rom_rdata <= 32'h00000000;
          16'h1c41 : blkif.rom_rdata <= 32'h00000000;
          16'h1c42 : blkif.rom_rdata <= 32'h00000000;
          16'h1c43 : blkif.rom_rdata <= 32'h00000000;
          16'h1c44 : blkif.rom_rdata <= 32'h00000000;
          16'h1c45 : blkif.rom_rdata <= 32'h00000000;
          16'h1c46 : blkif.rom_rdata <= 32'h00000000;
          16'h1c47 : blkif.rom_rdata <= 32'h00000000;
          16'h1c48 : blkif.rom_rdata <= 32'h00000000;
          16'h1c49 : blkif.rom_rdata <= 32'h00000000;
          16'h1c4a : blkif.rom_rdata <= 32'h00000000;
          16'h1c4b : blkif.rom_rdata <= 32'h00000000;
          16'h1c4c : blkif.rom_rdata <= 32'h00000000;
          16'h1c4d : blkif.rom_rdata <= 32'h00000000;
          16'h1c4e : blkif.rom_rdata <= 32'h00000000;
          16'h1c4f : blkif.rom_rdata <= 32'h00000000;
          16'h1c50 : blkif.rom_rdata <= 32'h00000000;
          16'h1c51 : blkif.rom_rdata <= 32'h00000000;
          16'h1c52 : blkif.rom_rdata <= 32'h00000000;
          16'h1c53 : blkif.rom_rdata <= 32'h00000000;
          16'h1c54 : blkif.rom_rdata <= 32'h00000000;
          16'h1c55 : blkif.rom_rdata <= 32'h00000000;
          16'h1c56 : blkif.rom_rdata <= 32'h00000000;
          16'h1c57 : blkif.rom_rdata <= 32'h00000000;
          16'h1c58 : blkif.rom_rdata <= 32'h00000000;
          16'h1c59 : blkif.rom_rdata <= 32'h00000000;
          16'h1c5a : blkif.rom_rdata <= 32'h00000000;
          16'h1c5b : blkif.rom_rdata <= 32'h00000000;
          16'h1c5c : blkif.rom_rdata <= 32'h00000000;
          16'h1c5d : blkif.rom_rdata <= 32'h00000000;
          16'h1c5e : blkif.rom_rdata <= 32'h00000000;
          16'h1c5f : blkif.rom_rdata <= 32'h00000000;
          16'h1c60 : blkif.rom_rdata <= 32'h00000000;
          16'h1c61 : blkif.rom_rdata <= 32'h00000000;
          16'h1c62 : blkif.rom_rdata <= 32'h00000000;
          16'h1c63 : blkif.rom_rdata <= 32'h00000000;
          16'h1c64 : blkif.rom_rdata <= 32'h00000000;
          16'h1c65 : blkif.rom_rdata <= 32'h00000000;
          16'h1c66 : blkif.rom_rdata <= 32'h00000000;
          16'h1c67 : blkif.rom_rdata <= 32'h00000000;
          16'h1c68 : blkif.rom_rdata <= 32'h00000000;
          16'h1c69 : blkif.rom_rdata <= 32'h00000000;
          16'h1c6a : blkif.rom_rdata <= 32'h00000000;
          16'h1c6b : blkif.rom_rdata <= 32'h00000000;
          16'h1c6c : blkif.rom_rdata <= 32'h00000000;
          16'h1c6d : blkif.rom_rdata <= 32'h00000000;
          16'h1c6e : blkif.rom_rdata <= 32'h00000000;
          16'h1c6f : blkif.rom_rdata <= 32'h00000000;
          16'h1c70 : blkif.rom_rdata <= 32'h00000000;
          16'h1c71 : blkif.rom_rdata <= 32'h00000000;
          16'h1c72 : blkif.rom_rdata <= 32'h00000000;
          16'h1c73 : blkif.rom_rdata <= 32'h00000000;
          16'h1c74 : blkif.rom_rdata <= 32'h00000000;
          16'h1c75 : blkif.rom_rdata <= 32'h00000000;
          16'h1c76 : blkif.rom_rdata <= 32'h00000000;
          16'h1c77 : blkif.rom_rdata <= 32'h00000000;
          16'h1c78 : blkif.rom_rdata <= 32'h00000000;
          16'h1c79 : blkif.rom_rdata <= 32'h00000000;
          16'h1c7a : blkif.rom_rdata <= 32'h00000000;
          16'h1c7b : blkif.rom_rdata <= 32'h00000000;
          16'h1c7c : blkif.rom_rdata <= 32'h00000000;
          16'h1c7d : blkif.rom_rdata <= 32'h00000000;
          16'h1c7e : blkif.rom_rdata <= 32'h00000000;
          16'h1c7f : blkif.rom_rdata <= 32'h00000000;
          16'h1c80 : blkif.rom_rdata <= 32'h00000000;
          16'h1c81 : blkif.rom_rdata <= 32'h00000000;
          16'h1c82 : blkif.rom_rdata <= 32'h00000000;
          16'h1c83 : blkif.rom_rdata <= 32'h00000000;
          16'h1c84 : blkif.rom_rdata <= 32'h00000000;
          16'h1c85 : blkif.rom_rdata <= 32'h00000000;
          16'h1c86 : blkif.rom_rdata <= 32'h00000000;
          16'h1c87 : blkif.rom_rdata <= 32'h00000000;
          16'h1c88 : blkif.rom_rdata <= 32'h00000000;
          16'h1c89 : blkif.rom_rdata <= 32'h00000000;
          16'h1c8a : blkif.rom_rdata <= 32'h00000000;
          16'h1c8b : blkif.rom_rdata <= 32'h00000000;
          16'h1c8c : blkif.rom_rdata <= 32'h00000000;
          16'h1c8d : blkif.rom_rdata <= 32'h00000000;
          16'h1c8e : blkif.rom_rdata <= 32'h00000000;
          16'h1c8f : blkif.rom_rdata <= 32'h00000000;
          16'h1c90 : blkif.rom_rdata <= 32'h00000000;
          16'h1c91 : blkif.rom_rdata <= 32'h00000000;
          16'h1c92 : blkif.rom_rdata <= 32'h00000000;
          16'h1c93 : blkif.rom_rdata <= 32'h00000000;
          16'h1c94 : blkif.rom_rdata <= 32'h00000000;
          16'h1c95 : blkif.rom_rdata <= 32'h00000000;
          16'h1c96 : blkif.rom_rdata <= 32'h00000000;
          16'h1c97 : blkif.rom_rdata <= 32'h00000000;
          16'h1c98 : blkif.rom_rdata <= 32'h00000000;
          16'h1c99 : blkif.rom_rdata <= 32'h00000000;
          16'h1c9a : blkif.rom_rdata <= 32'h00000000;
          16'h1c9b : blkif.rom_rdata <= 32'h00000000;
          16'h1c9c : blkif.rom_rdata <= 32'h00000000;
          16'h1c9d : blkif.rom_rdata <= 32'h00000000;
          16'h1c9e : blkif.rom_rdata <= 32'h00000000;
          16'h1c9f : blkif.rom_rdata <= 32'h00000000;
          16'h1ca0 : blkif.rom_rdata <= 32'h00000000;
          16'h1ca1 : blkif.rom_rdata <= 32'h00000000;
          16'h1ca2 : blkif.rom_rdata <= 32'h00000000;
          16'h1ca3 : blkif.rom_rdata <= 32'h00000000;
          16'h1ca4 : blkif.rom_rdata <= 32'h00000000;
          16'h1ca5 : blkif.rom_rdata <= 32'h00000000;
          16'h1ca6 : blkif.rom_rdata <= 32'h00000000;
          16'h1ca7 : blkif.rom_rdata <= 32'h00000000;
          16'h1ca8 : blkif.rom_rdata <= 32'h00000000;
          16'h1ca9 : blkif.rom_rdata <= 32'h00000000;
          16'h1caa : blkif.rom_rdata <= 32'h00000000;
          16'h1cab : blkif.rom_rdata <= 32'h00000000;
          16'h1cac : blkif.rom_rdata <= 32'h00000000;
          16'h1cad : blkif.rom_rdata <= 32'h00000000;
          16'h1cae : blkif.rom_rdata <= 32'h00000000;
          16'h1caf : blkif.rom_rdata <= 32'h00000000;
          16'h1cb0 : blkif.rom_rdata <= 32'h00000000;
          16'h1cb1 : blkif.rom_rdata <= 32'h00000000;
          16'h1cb2 : blkif.rom_rdata <= 32'h00000000;
          16'h1cb3 : blkif.rom_rdata <= 32'h00000000;
          16'h1cb4 : blkif.rom_rdata <= 32'h00000000;
          16'h1cb5 : blkif.rom_rdata <= 32'h00000000;
          16'h1cb6 : blkif.rom_rdata <= 32'h00000000;
          16'h1cb7 : blkif.rom_rdata <= 32'h00000000;
          16'h1cb8 : blkif.rom_rdata <= 32'h00000000;
          16'h1cb9 : blkif.rom_rdata <= 32'h00000000;
          16'h1cba : blkif.rom_rdata <= 32'h00000000;
          16'h1cbb : blkif.rom_rdata <= 32'h00000000;
          16'h1cbc : blkif.rom_rdata <= 32'h00000000;
          16'h1cbd : blkif.rom_rdata <= 32'h00000000;
          16'h1cbe : blkif.rom_rdata <= 32'h00000000;
          16'h1cbf : blkif.rom_rdata <= 32'h00000000;
          16'h1cc0 : blkif.rom_rdata <= 32'h00000000;
          16'h1cc1 : blkif.rom_rdata <= 32'h00000000;
          16'h1cc2 : blkif.rom_rdata <= 32'h00000000;
          16'h1cc3 : blkif.rom_rdata <= 32'h00000000;
          16'h1cc4 : blkif.rom_rdata <= 32'h00000000;
          16'h1cc5 : blkif.rom_rdata <= 32'h00000000;
          16'h1cc6 : blkif.rom_rdata <= 32'h00000000;
          16'h1cc7 : blkif.rom_rdata <= 32'h00000000;
          16'h1cc8 : blkif.rom_rdata <= 32'h00000000;
          16'h1cc9 : blkif.rom_rdata <= 32'h00000000;
          16'h1cca : blkif.rom_rdata <= 32'h00000000;
          16'h1ccb : blkif.rom_rdata <= 32'h00000000;
          16'h1ccc : blkif.rom_rdata <= 32'h00000000;
          16'h1ccd : blkif.rom_rdata <= 32'h00000000;
          16'h1cce : blkif.rom_rdata <= 32'h00000000;
          16'h1ccf : blkif.rom_rdata <= 32'h00000000;
          16'h1cd0 : blkif.rom_rdata <= 32'h00000000;
          16'h1cd1 : blkif.rom_rdata <= 32'h00000000;
          16'h1cd2 : blkif.rom_rdata <= 32'h00000000;
          16'h1cd3 : blkif.rom_rdata <= 32'h00000000;
          16'h1cd4 : blkif.rom_rdata <= 32'h00000000;
          16'h1cd5 : blkif.rom_rdata <= 32'h00000000;
          16'h1cd6 : blkif.rom_rdata <= 32'h00000000;
          16'h1cd7 : blkif.rom_rdata <= 32'h00000000;
          16'h1cd8 : blkif.rom_rdata <= 32'h00000000;
          16'h1cd9 : blkif.rom_rdata <= 32'h00000000;
          16'h1cda : blkif.rom_rdata <= 32'h00000000;
          16'h1cdb : blkif.rom_rdata <= 32'h00000000;
          16'h1cdc : blkif.rom_rdata <= 32'h00000000;
          16'h1cdd : blkif.rom_rdata <= 32'h00000000;
          16'h1cde : blkif.rom_rdata <= 32'h00000000;
          16'h1cdf : blkif.rom_rdata <= 32'h00000000;
          16'h1ce0 : blkif.rom_rdata <= 32'h00000000;
          16'h1ce1 : blkif.rom_rdata <= 32'h00000000;
          16'h1ce2 : blkif.rom_rdata <= 32'h00000000;
          16'h1ce3 : blkif.rom_rdata <= 32'h00000000;
          16'h1ce4 : blkif.rom_rdata <= 32'h00000000;
          16'h1ce5 : blkif.rom_rdata <= 32'h00000000;
          16'h1ce6 : blkif.rom_rdata <= 32'h00000000;
          16'h1ce7 : blkif.rom_rdata <= 32'h00000000;
          16'h1ce8 : blkif.rom_rdata <= 32'h00000000;
          16'h1ce9 : blkif.rom_rdata <= 32'h00000000;
          16'h1cea : blkif.rom_rdata <= 32'h00000000;
          16'h1ceb : blkif.rom_rdata <= 32'h00000000;
          16'h1cec : blkif.rom_rdata <= 32'h00000000;
          16'h1ced : blkif.rom_rdata <= 32'h00000000;
          16'h1cee : blkif.rom_rdata <= 32'h00000000;
          16'h1cef : blkif.rom_rdata <= 32'h00000000;
          16'h1cf0 : blkif.rom_rdata <= 32'h00000000;
          16'h1cf1 : blkif.rom_rdata <= 32'h00000000;
          16'h1cf2 : blkif.rom_rdata <= 32'h00000000;
          16'h1cf3 : blkif.rom_rdata <= 32'h00000000;
          16'h1cf4 : blkif.rom_rdata <= 32'h00000000;
          16'h1cf5 : blkif.rom_rdata <= 32'h00000000;
          16'h1cf6 : blkif.rom_rdata <= 32'h00000000;
          16'h1cf7 : blkif.rom_rdata <= 32'h00000000;
          16'h1cf8 : blkif.rom_rdata <= 32'h00000000;
          16'h1cf9 : blkif.rom_rdata <= 32'h00000000;
          16'h1cfa : blkif.rom_rdata <= 32'h00000000;
          16'h1cfb : blkif.rom_rdata <= 32'h00000000;
          16'h1cfc : blkif.rom_rdata <= 32'h00000000;
          16'h1cfd : blkif.rom_rdata <= 32'h00000000;
          16'h1cfe : blkif.rom_rdata <= 32'h00000000;
          16'h1cff : blkif.rom_rdata <= 32'h00000000;
          16'h1d00 : blkif.rom_rdata <= 32'h00000000;
          16'h1d01 : blkif.rom_rdata <= 32'h00000000;
          16'h1d02 : blkif.rom_rdata <= 32'h00000000;
          16'h1d03 : blkif.rom_rdata <= 32'h00000000;
          16'h1d04 : blkif.rom_rdata <= 32'h00000000;
          16'h1d05 : blkif.rom_rdata <= 32'h00000000;
          16'h1d06 : blkif.rom_rdata <= 32'h00000000;
          16'h1d07 : blkif.rom_rdata <= 32'h00000000;
          16'h1d08 : blkif.rom_rdata <= 32'h00000000;
          16'h1d09 : blkif.rom_rdata <= 32'h00000000;
          16'h1d0a : blkif.rom_rdata <= 32'h00000000;
          16'h1d0b : blkif.rom_rdata <= 32'h00000000;
          16'h1d0c : blkif.rom_rdata <= 32'h00000000;
          16'h1d0d : blkif.rom_rdata <= 32'h00000000;
          16'h1d0e : blkif.rom_rdata <= 32'h00000000;
          16'h1d0f : blkif.rom_rdata <= 32'h00000000;
          16'h1d10 : blkif.rom_rdata <= 32'h00000000;
          16'h1d11 : blkif.rom_rdata <= 32'h00000000;
          16'h1d12 : blkif.rom_rdata <= 32'h00000000;
          16'h1d13 : blkif.rom_rdata <= 32'h00000000;
          16'h1d14 : blkif.rom_rdata <= 32'h00000000;
          16'h1d15 : blkif.rom_rdata <= 32'h00000000;
          16'h1d16 : blkif.rom_rdata <= 32'h00000000;
          16'h1d17 : blkif.rom_rdata <= 32'h00000000;
          16'h1d18 : blkif.rom_rdata <= 32'h00000000;
          16'h1d19 : blkif.rom_rdata <= 32'h00000000;
          16'h1d1a : blkif.rom_rdata <= 32'h00000000;
          16'h1d1b : blkif.rom_rdata <= 32'h00000000;
          16'h1d1c : blkif.rom_rdata <= 32'h00000000;
          16'h1d1d : blkif.rom_rdata <= 32'h00000000;
          16'h1d1e : blkif.rom_rdata <= 32'h00000000;
          16'h1d1f : blkif.rom_rdata <= 32'h00000000;
          16'h1d20 : blkif.rom_rdata <= 32'h00000000;
          16'h1d21 : blkif.rom_rdata <= 32'h00000000;
          16'h1d22 : blkif.rom_rdata <= 32'h00000000;
          16'h1d23 : blkif.rom_rdata <= 32'h00000000;
          16'h1d24 : blkif.rom_rdata <= 32'h00000000;
          16'h1d25 : blkif.rom_rdata <= 32'h00000000;
          16'h1d26 : blkif.rom_rdata <= 32'h00000000;
          16'h1d27 : blkif.rom_rdata <= 32'h00000000;
          16'h1d28 : blkif.rom_rdata <= 32'h00000000;
          16'h1d29 : blkif.rom_rdata <= 32'h00000000;
          16'h1d2a : blkif.rom_rdata <= 32'h00000000;
          16'h1d2b : blkif.rom_rdata <= 32'h00000000;
          16'h1d2c : blkif.rom_rdata <= 32'h00000000;
          16'h1d2d : blkif.rom_rdata <= 32'h00000000;
          16'h1d2e : blkif.rom_rdata <= 32'h00000000;
          16'h1d2f : blkif.rom_rdata <= 32'h00000000;
          16'h1d30 : blkif.rom_rdata <= 32'h00000000;
          16'h1d31 : blkif.rom_rdata <= 32'h00000000;
          16'h1d32 : blkif.rom_rdata <= 32'h00000000;
          16'h1d33 : blkif.rom_rdata <= 32'h00000000;
          16'h1d34 : blkif.rom_rdata <= 32'h00000000;
          16'h1d35 : blkif.rom_rdata <= 32'h00000000;
          16'h1d36 : blkif.rom_rdata <= 32'h00000000;
          16'h1d37 : blkif.rom_rdata <= 32'h00000000;
          16'h1d38 : blkif.rom_rdata <= 32'h00000000;
          16'h1d39 : blkif.rom_rdata <= 32'h00000000;
          16'h1d3a : blkif.rom_rdata <= 32'h00000000;
          16'h1d3b : blkif.rom_rdata <= 32'h00000000;
          16'h1d3c : blkif.rom_rdata <= 32'h00000000;
          16'h1d3d : blkif.rom_rdata <= 32'h00000000;
          16'h1d3e : blkif.rom_rdata <= 32'h00000000;
          16'h1d3f : blkif.rom_rdata <= 32'h00000000;
          16'h1d40 : blkif.rom_rdata <= 32'h00000000;
          16'h1d41 : blkif.rom_rdata <= 32'h00000000;
          16'h1d42 : blkif.rom_rdata <= 32'h00000000;
          16'h1d43 : blkif.rom_rdata <= 32'h00000000;
          16'h1d44 : blkif.rom_rdata <= 32'h00000000;
          16'h1d45 : blkif.rom_rdata <= 32'h00000000;
          16'h1d46 : blkif.rom_rdata <= 32'h00000000;
          16'h1d47 : blkif.rom_rdata <= 32'h00000000;
          16'h1d48 : blkif.rom_rdata <= 32'h00000000;
          16'h1d49 : blkif.rom_rdata <= 32'h00000000;
          16'h1d4a : blkif.rom_rdata <= 32'h00000000;
          16'h1d4b : blkif.rom_rdata <= 32'h00000000;
          16'h1d4c : blkif.rom_rdata <= 32'h00000000;
          16'h1d4d : blkif.rom_rdata <= 32'h00000000;
          16'h1d4e : blkif.rom_rdata <= 32'h00000000;
          16'h1d4f : blkif.rom_rdata <= 32'h00000000;
          16'h1d50 : blkif.rom_rdata <= 32'h00000000;
          16'h1d51 : blkif.rom_rdata <= 32'h00000000;
          16'h1d52 : blkif.rom_rdata <= 32'h00000000;
          16'h1d53 : blkif.rom_rdata <= 32'h00000000;
          16'h1d54 : blkif.rom_rdata <= 32'h00000000;
          16'h1d55 : blkif.rom_rdata <= 32'h00000000;
          16'h1d56 : blkif.rom_rdata <= 32'h00000000;
          16'h1d57 : blkif.rom_rdata <= 32'h00000000;
          16'h1d58 : blkif.rom_rdata <= 32'h00000000;
          16'h1d59 : blkif.rom_rdata <= 32'h00000000;
          16'h1d5a : blkif.rom_rdata <= 32'h00000000;
          16'h1d5b : blkif.rom_rdata <= 32'h00000000;
          16'h1d5c : blkif.rom_rdata <= 32'h00000000;
          16'h1d5d : blkif.rom_rdata <= 32'h00000000;
          16'h1d5e : blkif.rom_rdata <= 32'h00000000;
          16'h1d5f : blkif.rom_rdata <= 32'h00000000;
          16'h1d60 : blkif.rom_rdata <= 32'h00000000;
          16'h1d61 : blkif.rom_rdata <= 32'h00000000;
          16'h1d62 : blkif.rom_rdata <= 32'h00000000;
          16'h1d63 : blkif.rom_rdata <= 32'h00000000;
          16'h1d64 : blkif.rom_rdata <= 32'h00000000;
          16'h1d65 : blkif.rom_rdata <= 32'h00000000;
          16'h1d66 : blkif.rom_rdata <= 32'h00000000;
          16'h1d67 : blkif.rom_rdata <= 32'h00000000;
          16'h1d68 : blkif.rom_rdata <= 32'h00000000;
          16'h1d69 : blkif.rom_rdata <= 32'h00000000;
          16'h1d6a : blkif.rom_rdata <= 32'h00000000;
          16'h1d6b : blkif.rom_rdata <= 32'h00000000;
          16'h1d6c : blkif.rom_rdata <= 32'h00000000;
          16'h1d6d : blkif.rom_rdata <= 32'h00000000;
          16'h1d6e : blkif.rom_rdata <= 32'h00000000;
          16'h1d6f : blkif.rom_rdata <= 32'h00000000;
          16'h1d70 : blkif.rom_rdata <= 32'h00000000;
          16'h1d71 : blkif.rom_rdata <= 32'h00000000;
          16'h1d72 : blkif.rom_rdata <= 32'h00000000;
          16'h1d73 : blkif.rom_rdata <= 32'h00000000;
          16'h1d74 : blkif.rom_rdata <= 32'h00000000;
          16'h1d75 : blkif.rom_rdata <= 32'h00000000;
          16'h1d76 : blkif.rom_rdata <= 32'h00000000;
          16'h1d77 : blkif.rom_rdata <= 32'h00000000;
          16'h1d78 : blkif.rom_rdata <= 32'h00000000;
          16'h1d79 : blkif.rom_rdata <= 32'h00000000;
          16'h1d7a : blkif.rom_rdata <= 32'h00000000;
          16'h1d7b : blkif.rom_rdata <= 32'h00000000;
          16'h1d7c : blkif.rom_rdata <= 32'h00000000;
          16'h1d7d : blkif.rom_rdata <= 32'h00000000;
          16'h1d7e : blkif.rom_rdata <= 32'h00000000;
          16'h1d7f : blkif.rom_rdata <= 32'h00000000;
          16'h1d80 : blkif.rom_rdata <= 32'h00000000;
          16'h1d81 : blkif.rom_rdata <= 32'h00000000;
          16'h1d82 : blkif.rom_rdata <= 32'h00000000;
          16'h1d83 : blkif.rom_rdata <= 32'h00000000;
          16'h1d84 : blkif.rom_rdata <= 32'h00000000;
          16'h1d85 : blkif.rom_rdata <= 32'h00000000;
          16'h1d86 : blkif.rom_rdata <= 32'h00000000;
          16'h1d87 : blkif.rom_rdata <= 32'h00000000;
          16'h1d88 : blkif.rom_rdata <= 32'h00000000;
          16'h1d89 : blkif.rom_rdata <= 32'h00000000;
          16'h1d8a : blkif.rom_rdata <= 32'h00000000;
          16'h1d8b : blkif.rom_rdata <= 32'h00000000;
          16'h1d8c : blkif.rom_rdata <= 32'h00000000;
          16'h1d8d : blkif.rom_rdata <= 32'h00000000;
          16'h1d8e : blkif.rom_rdata <= 32'h00000000;
          16'h1d8f : blkif.rom_rdata <= 32'h00000000;
          16'h1d90 : blkif.rom_rdata <= 32'h00000000;
          16'h1d91 : blkif.rom_rdata <= 32'h00000000;
          16'h1d92 : blkif.rom_rdata <= 32'h00000000;
          16'h1d93 : blkif.rom_rdata <= 32'h00000000;
          16'h1d94 : blkif.rom_rdata <= 32'h00000000;
          16'h1d95 : blkif.rom_rdata <= 32'h00000000;
          16'h1d96 : blkif.rom_rdata <= 32'h00000000;
          16'h1d97 : blkif.rom_rdata <= 32'h00000000;
          16'h1d98 : blkif.rom_rdata <= 32'h00000000;
          16'h1d99 : blkif.rom_rdata <= 32'h00000000;
          16'h1d9a : blkif.rom_rdata <= 32'h00000000;
          16'h1d9b : blkif.rom_rdata <= 32'h00000000;
          16'h1d9c : blkif.rom_rdata <= 32'h00000000;
          16'h1d9d : blkif.rom_rdata <= 32'h00000000;
          16'h1d9e : blkif.rom_rdata <= 32'h00000000;
          16'h1d9f : blkif.rom_rdata <= 32'h00000000;
          16'h1da0 : blkif.rom_rdata <= 32'h00000000;
          16'h1da1 : blkif.rom_rdata <= 32'h00000000;
          16'h1da2 : blkif.rom_rdata <= 32'h00000000;
          16'h1da3 : blkif.rom_rdata <= 32'h00000000;
          16'h1da4 : blkif.rom_rdata <= 32'h00000000;
          16'h1da5 : blkif.rom_rdata <= 32'h00000000;
          16'h1da6 : blkif.rom_rdata <= 32'h00000000;
          16'h1da7 : blkif.rom_rdata <= 32'h00000000;
          16'h1da8 : blkif.rom_rdata <= 32'h00000000;
          16'h1da9 : blkif.rom_rdata <= 32'h00000000;
          16'h1daa : blkif.rom_rdata <= 32'h00000000;
          16'h1dab : blkif.rom_rdata <= 32'h00000000;
          16'h1dac : blkif.rom_rdata <= 32'h00000000;
          16'h1dad : blkif.rom_rdata <= 32'h00000000;
          16'h1dae : blkif.rom_rdata <= 32'h00000000;
          16'h1daf : blkif.rom_rdata <= 32'h00000000;
          16'h1db0 : blkif.rom_rdata <= 32'h00000000;
          16'h1db1 : blkif.rom_rdata <= 32'h00000000;
          16'h1db2 : blkif.rom_rdata <= 32'h00000000;
          16'h1db3 : blkif.rom_rdata <= 32'h00000000;
          16'h1db4 : blkif.rom_rdata <= 32'h00000000;
          16'h1db5 : blkif.rom_rdata <= 32'h00000000;
          16'h1db6 : blkif.rom_rdata <= 32'h00000000;
          16'h1db7 : blkif.rom_rdata <= 32'h00000000;
          16'h1db8 : blkif.rom_rdata <= 32'h00000000;
          16'h1db9 : blkif.rom_rdata <= 32'h00000000;
          16'h1dba : blkif.rom_rdata <= 32'h00000000;
          16'h1dbb : blkif.rom_rdata <= 32'h00000000;
          16'h1dbc : blkif.rom_rdata <= 32'h00000000;
          16'h1dbd : blkif.rom_rdata <= 32'h00000000;
          16'h1dbe : blkif.rom_rdata <= 32'h00000000;
          16'h1dbf : blkif.rom_rdata <= 32'h00000000;
          16'h1dc0 : blkif.rom_rdata <= 32'h00000000;
          16'h1dc1 : blkif.rom_rdata <= 32'h00000000;
          16'h1dc2 : blkif.rom_rdata <= 32'h00000000;
          16'h1dc3 : blkif.rom_rdata <= 32'h00000000;
          16'h1dc4 : blkif.rom_rdata <= 32'h00000000;
          16'h1dc5 : blkif.rom_rdata <= 32'h00000000;
          16'h1dc6 : blkif.rom_rdata <= 32'h00000000;
          16'h1dc7 : blkif.rom_rdata <= 32'h00000000;
          16'h1dc8 : blkif.rom_rdata <= 32'h00000000;
          16'h1dc9 : blkif.rom_rdata <= 32'h00000000;
          16'h1dca : blkif.rom_rdata <= 32'h00000000;
          16'h1dcb : blkif.rom_rdata <= 32'h00000000;
          16'h1dcc : blkif.rom_rdata <= 32'h00000000;
          16'h1dcd : blkif.rom_rdata <= 32'h00000000;
          16'h1dce : blkif.rom_rdata <= 32'h00000000;
          16'h1dcf : blkif.rom_rdata <= 32'h00000000;
          16'h1dd0 : blkif.rom_rdata <= 32'h00000000;
          16'h1dd1 : blkif.rom_rdata <= 32'h00000000;
          16'h1dd2 : blkif.rom_rdata <= 32'h00000000;
          16'h1dd3 : blkif.rom_rdata <= 32'h00000000;
          16'h1dd4 : blkif.rom_rdata <= 32'h00000000;
          16'h1dd5 : blkif.rom_rdata <= 32'h00000000;
          16'h1dd6 : blkif.rom_rdata <= 32'h00000000;
          16'h1dd7 : blkif.rom_rdata <= 32'h00000000;
          16'h1dd8 : blkif.rom_rdata <= 32'h00000000;
          16'h1dd9 : blkif.rom_rdata <= 32'h00000000;
          16'h1dda : blkif.rom_rdata <= 32'h00000000;
          16'h1ddb : blkif.rom_rdata <= 32'h00000000;
          16'h1ddc : blkif.rom_rdata <= 32'h00000000;
          16'h1ddd : blkif.rom_rdata <= 32'h00000000;
          16'h1dde : blkif.rom_rdata <= 32'h00000000;
          16'h1ddf : blkif.rom_rdata <= 32'h00000000;
          16'h1de0 : blkif.rom_rdata <= 32'h00000000;
          16'h1de1 : blkif.rom_rdata <= 32'h00000000;
          16'h1de2 : blkif.rom_rdata <= 32'h00000000;
          16'h1de3 : blkif.rom_rdata <= 32'h00000000;
          16'h1de4 : blkif.rom_rdata <= 32'h00000000;
          16'h1de5 : blkif.rom_rdata <= 32'h00000000;
          16'h1de6 : blkif.rom_rdata <= 32'h00000000;
          16'h1de7 : blkif.rom_rdata <= 32'h00000000;
          16'h1de8 : blkif.rom_rdata <= 32'h00000000;
          16'h1de9 : blkif.rom_rdata <= 32'h00000000;
          16'h1dea : blkif.rom_rdata <= 32'h00000000;
          16'h1deb : blkif.rom_rdata <= 32'h00000000;
          16'h1dec : blkif.rom_rdata <= 32'h00000000;
          16'h1ded : blkif.rom_rdata <= 32'h00000000;
          16'h1dee : blkif.rom_rdata <= 32'h00000000;
          16'h1def : blkif.rom_rdata <= 32'h00000000;
          16'h1df0 : blkif.rom_rdata <= 32'h00000000;
          16'h1df1 : blkif.rom_rdata <= 32'h00000000;
          16'h1df2 : blkif.rom_rdata <= 32'h00000000;
          16'h1df3 : blkif.rom_rdata <= 32'h00000000;
          16'h1df4 : blkif.rom_rdata <= 32'h00000000;
          16'h1df5 : blkif.rom_rdata <= 32'h00000000;
          16'h1df6 : blkif.rom_rdata <= 32'h00000000;
          16'h1df7 : blkif.rom_rdata <= 32'h00000000;
          16'h1df8 : blkif.rom_rdata <= 32'h00000000;
          16'h1df9 : blkif.rom_rdata <= 32'h00000000;
          16'h1dfa : blkif.rom_rdata <= 32'h00000000;
          16'h1dfb : blkif.rom_rdata <= 32'h00000000;
          16'h1dfc : blkif.rom_rdata <= 32'h00000000;
          16'h1dfd : blkif.rom_rdata <= 32'h00000000;
          16'h1dfe : blkif.rom_rdata <= 32'h00000000;
          16'h1dff : blkif.rom_rdata <= 32'h00000000;
          16'h1e00 : blkif.rom_rdata <= 32'h00000000;
          16'h1e01 : blkif.rom_rdata <= 32'h00000000;
          16'h1e02 : blkif.rom_rdata <= 32'h00000000;
          16'h1e03 : blkif.rom_rdata <= 32'h00000000;
          16'h1e04 : blkif.rom_rdata <= 32'h00000000;
          16'h1e05 : blkif.rom_rdata <= 32'h00000000;
          16'h1e06 : blkif.rom_rdata <= 32'h00000000;
          16'h1e07 : blkif.rom_rdata <= 32'h00000000;
          16'h1e08 : blkif.rom_rdata <= 32'h00000000;
          16'h1e09 : blkif.rom_rdata <= 32'h00000000;
          16'h1e0a : blkif.rom_rdata <= 32'h00000000;
          16'h1e0b : blkif.rom_rdata <= 32'h00000000;
          16'h1e0c : blkif.rom_rdata <= 32'h00000000;
          16'h1e0d : blkif.rom_rdata <= 32'h00000000;
          16'h1e0e : blkif.rom_rdata <= 32'h00000000;
          16'h1e0f : blkif.rom_rdata <= 32'h00000000;
          16'h1e10 : blkif.rom_rdata <= 32'h00000000;
          16'h1e11 : blkif.rom_rdata <= 32'h00000000;
          16'h1e12 : blkif.rom_rdata <= 32'h00000000;
          16'h1e13 : blkif.rom_rdata <= 32'h00000000;
          16'h1e14 : blkif.rom_rdata <= 32'h00000000;
          16'h1e15 : blkif.rom_rdata <= 32'h00000000;
          16'h1e16 : blkif.rom_rdata <= 32'h00000000;
          16'h1e17 : blkif.rom_rdata <= 32'h00000000;
          16'h1e18 : blkif.rom_rdata <= 32'h00000000;
          16'h1e19 : blkif.rom_rdata <= 32'h00000000;
          16'h1e1a : blkif.rom_rdata <= 32'h00000000;
          16'h1e1b : blkif.rom_rdata <= 32'h00000000;
          16'h1e1c : blkif.rom_rdata <= 32'h00000000;
          16'h1e1d : blkif.rom_rdata <= 32'h00000000;
          16'h1e1e : blkif.rom_rdata <= 32'h00000000;
          16'h1e1f : blkif.rom_rdata <= 32'h00000000;
          16'h1e20 : blkif.rom_rdata <= 32'h00000000;
          16'h1e21 : blkif.rom_rdata <= 32'h00000000;
          16'h1e22 : blkif.rom_rdata <= 32'h00000000;
          16'h1e23 : blkif.rom_rdata <= 32'h00000000;
          16'h1e24 : blkif.rom_rdata <= 32'h00000000;
          16'h1e25 : blkif.rom_rdata <= 32'h00000000;
          16'h1e26 : blkif.rom_rdata <= 32'h00000000;
          16'h1e27 : blkif.rom_rdata <= 32'h00000000;
          16'h1e28 : blkif.rom_rdata <= 32'h00000000;
          16'h1e29 : blkif.rom_rdata <= 32'h00000000;
          16'h1e2a : blkif.rom_rdata <= 32'h00000000;
          16'h1e2b : blkif.rom_rdata <= 32'h00000000;
          16'h1e2c : blkif.rom_rdata <= 32'h00000000;
          16'h1e2d : blkif.rom_rdata <= 32'h00000000;
          16'h1e2e : blkif.rom_rdata <= 32'h00000000;
          16'h1e2f : blkif.rom_rdata <= 32'h00000000;
          16'h1e30 : blkif.rom_rdata <= 32'h00000000;
          16'h1e31 : blkif.rom_rdata <= 32'h00000000;
          16'h1e32 : blkif.rom_rdata <= 32'h00000000;
          16'h1e33 : blkif.rom_rdata <= 32'h00000000;
          16'h1e34 : blkif.rom_rdata <= 32'h00000000;
          16'h1e35 : blkif.rom_rdata <= 32'h00000000;
          16'h1e36 : blkif.rom_rdata <= 32'h00000000;
          16'h1e37 : blkif.rom_rdata <= 32'h00000000;
          16'h1e38 : blkif.rom_rdata <= 32'h00000000;
          16'h1e39 : blkif.rom_rdata <= 32'h00000000;
          16'h1e3a : blkif.rom_rdata <= 32'h00000000;
          16'h1e3b : blkif.rom_rdata <= 32'h00000000;
          16'h1e3c : blkif.rom_rdata <= 32'h00000000;
          16'h1e3d : blkif.rom_rdata <= 32'h00000000;
          16'h1e3e : blkif.rom_rdata <= 32'h00000000;
          16'h1e3f : blkif.rom_rdata <= 32'h00000000;
          16'h1e40 : blkif.rom_rdata <= 32'h00000000;
          16'h1e41 : blkif.rom_rdata <= 32'h00000000;
          16'h1e42 : blkif.rom_rdata <= 32'h00000000;
          16'h1e43 : blkif.rom_rdata <= 32'h00000000;
          16'h1e44 : blkif.rom_rdata <= 32'h00000000;
          16'h1e45 : blkif.rom_rdata <= 32'h00000000;
          16'h1e46 : blkif.rom_rdata <= 32'h00000000;
          16'h1e47 : blkif.rom_rdata <= 32'h00000000;
          16'h1e48 : blkif.rom_rdata <= 32'h00000000;
          16'h1e49 : blkif.rom_rdata <= 32'h00000000;
          16'h1e4a : blkif.rom_rdata <= 32'h00000000;
          16'h1e4b : blkif.rom_rdata <= 32'h00000000;
          16'h1e4c : blkif.rom_rdata <= 32'h00000000;
          16'h1e4d : blkif.rom_rdata <= 32'h00000000;
          16'h1e4e : blkif.rom_rdata <= 32'h00000000;
          16'h1e4f : blkif.rom_rdata <= 32'h00000000;
          16'h1e50 : blkif.rom_rdata <= 32'h00000000;
          16'h1e51 : blkif.rom_rdata <= 32'h00000000;
          16'h1e52 : blkif.rom_rdata <= 32'h00000000;
          16'h1e53 : blkif.rom_rdata <= 32'h00000000;
          16'h1e54 : blkif.rom_rdata <= 32'h00000000;
          16'h1e55 : blkif.rom_rdata <= 32'h00000000;
          16'h1e56 : blkif.rom_rdata <= 32'h00000000;
          16'h1e57 : blkif.rom_rdata <= 32'h00000000;
          16'h1e58 : blkif.rom_rdata <= 32'h00000000;
          16'h1e59 : blkif.rom_rdata <= 32'h00000000;
          16'h1e5a : blkif.rom_rdata <= 32'h00000000;
          16'h1e5b : blkif.rom_rdata <= 32'h00000000;
          16'h1e5c : blkif.rom_rdata <= 32'h00000000;
          16'h1e5d : blkif.rom_rdata <= 32'h00000000;
          16'h1e5e : blkif.rom_rdata <= 32'h00000000;
          16'h1e5f : blkif.rom_rdata <= 32'h00000000;
          16'h1e60 : blkif.rom_rdata <= 32'h00000000;
          16'h1e61 : blkif.rom_rdata <= 32'h00000000;
          16'h1e62 : blkif.rom_rdata <= 32'h00000000;
          16'h1e63 : blkif.rom_rdata <= 32'h00000000;
          16'h1e64 : blkif.rom_rdata <= 32'h00000000;
          16'h1e65 : blkif.rom_rdata <= 32'h00000000;
          16'h1e66 : blkif.rom_rdata <= 32'h00000000;
          16'h1e67 : blkif.rom_rdata <= 32'h00000000;
          16'h1e68 : blkif.rom_rdata <= 32'h00000000;
          16'h1e69 : blkif.rom_rdata <= 32'h00000000;
          16'h1e6a : blkif.rom_rdata <= 32'h00000000;
          16'h1e6b : blkif.rom_rdata <= 32'h00000000;
          16'h1e6c : blkif.rom_rdata <= 32'h00000000;
          16'h1e6d : blkif.rom_rdata <= 32'h00000000;
          16'h1e6e : blkif.rom_rdata <= 32'h00000000;
          16'h1e6f : blkif.rom_rdata <= 32'h00000000;
          16'h1e70 : blkif.rom_rdata <= 32'h00000000;
          16'h1e71 : blkif.rom_rdata <= 32'h00000000;
          16'h1e72 : blkif.rom_rdata <= 32'h00000000;
          16'h1e73 : blkif.rom_rdata <= 32'h00000000;
          16'h1e74 : blkif.rom_rdata <= 32'h00000000;
          16'h1e75 : blkif.rom_rdata <= 32'h00000000;
          16'h1e76 : blkif.rom_rdata <= 32'h00000000;
          16'h1e77 : blkif.rom_rdata <= 32'h00000000;
          16'h1e78 : blkif.rom_rdata <= 32'h00000000;
          16'h1e79 : blkif.rom_rdata <= 32'h00000000;
          16'h1e7a : blkif.rom_rdata <= 32'h00000000;
          16'h1e7b : blkif.rom_rdata <= 32'h00000000;
          16'h1e7c : blkif.rom_rdata <= 32'h00000000;
          16'h1e7d : blkif.rom_rdata <= 32'h00000000;
          16'h1e7e : blkif.rom_rdata <= 32'h00000000;
          16'h1e7f : blkif.rom_rdata <= 32'h00000000;
          16'h1e80 : blkif.rom_rdata <= 32'h00000000;
          16'h1e81 : blkif.rom_rdata <= 32'h00000000;
          16'h1e82 : blkif.rom_rdata <= 32'h00000000;
          16'h1e83 : blkif.rom_rdata <= 32'h00000000;
          16'h1e84 : blkif.rom_rdata <= 32'h00000000;
          16'h1e85 : blkif.rom_rdata <= 32'h00000000;
          16'h1e86 : blkif.rom_rdata <= 32'h00000000;
          16'h1e87 : blkif.rom_rdata <= 32'h00000000;
          16'h1e88 : blkif.rom_rdata <= 32'h00000000;
          16'h1e89 : blkif.rom_rdata <= 32'h00000000;
          16'h1e8a : blkif.rom_rdata <= 32'h00000000;
          16'h1e8b : blkif.rom_rdata <= 32'h00000000;
          16'h1e8c : blkif.rom_rdata <= 32'h00000000;
          16'h1e8d : blkif.rom_rdata <= 32'h00000000;
          16'h1e8e : blkif.rom_rdata <= 32'h00000000;
          16'h1e8f : blkif.rom_rdata <= 32'h00000000;
          16'h1e90 : blkif.rom_rdata <= 32'h00000000;
          16'h1e91 : blkif.rom_rdata <= 32'h00000000;
          16'h1e92 : blkif.rom_rdata <= 32'h00000000;
          16'h1e93 : blkif.rom_rdata <= 32'h00000000;
          16'h1e94 : blkif.rom_rdata <= 32'h00000000;
          16'h1e95 : blkif.rom_rdata <= 32'h00000000;
          16'h1e96 : blkif.rom_rdata <= 32'h00000000;
          16'h1e97 : blkif.rom_rdata <= 32'h00000000;
          16'h1e98 : blkif.rom_rdata <= 32'h00000000;
          16'h1e99 : blkif.rom_rdata <= 32'h00000000;
          16'h1e9a : blkif.rom_rdata <= 32'h00000000;
          16'h1e9b : blkif.rom_rdata <= 32'h00000000;
          16'h1e9c : blkif.rom_rdata <= 32'h00000000;
          16'h1e9d : blkif.rom_rdata <= 32'h00000000;
          16'h1e9e : blkif.rom_rdata <= 32'h00000000;
          16'h1e9f : blkif.rom_rdata <= 32'h00000000;
          16'h1ea0 : blkif.rom_rdata <= 32'h00000000;
          16'h1ea1 : blkif.rom_rdata <= 32'h00000000;
          16'h1ea2 : blkif.rom_rdata <= 32'h00000000;
          16'h1ea3 : blkif.rom_rdata <= 32'h00000000;
          16'h1ea4 : blkif.rom_rdata <= 32'h00000000;
          16'h1ea5 : blkif.rom_rdata <= 32'h00000000;
          16'h1ea6 : blkif.rom_rdata <= 32'h00000000;
          16'h1ea7 : blkif.rom_rdata <= 32'h00000000;
          16'h1ea8 : blkif.rom_rdata <= 32'h00000000;
          16'h1ea9 : blkif.rom_rdata <= 32'h00000000;
          16'h1eaa : blkif.rom_rdata <= 32'h00000000;
          16'h1eab : blkif.rom_rdata <= 32'h00000000;
          16'h1eac : blkif.rom_rdata <= 32'h00000000;
          16'h1ead : blkif.rom_rdata <= 32'h00000000;
          16'h1eae : blkif.rom_rdata <= 32'h00000000;
          16'h1eaf : blkif.rom_rdata <= 32'h00000000;
          16'h1eb0 : blkif.rom_rdata <= 32'h00000000;
          16'h1eb1 : blkif.rom_rdata <= 32'h00000000;
          16'h1eb2 : blkif.rom_rdata <= 32'h00000000;
          16'h1eb3 : blkif.rom_rdata <= 32'h00000000;
          16'h1eb4 : blkif.rom_rdata <= 32'h00000000;
          16'h1eb5 : blkif.rom_rdata <= 32'h00000000;
          16'h1eb6 : blkif.rom_rdata <= 32'h00000000;
          16'h1eb7 : blkif.rom_rdata <= 32'h00000000;
          16'h1eb8 : blkif.rom_rdata <= 32'h00000000;
          16'h1eb9 : blkif.rom_rdata <= 32'h00000000;
          16'h1eba : blkif.rom_rdata <= 32'h00000000;
          16'h1ebb : blkif.rom_rdata <= 32'h00000000;
          16'h1ebc : blkif.rom_rdata <= 32'h00000000;
          16'h1ebd : blkif.rom_rdata <= 32'h00000000;
          16'h1ebe : blkif.rom_rdata <= 32'h00000000;
          16'h1ebf : blkif.rom_rdata <= 32'h00000000;
          16'h1ec0 : blkif.rom_rdata <= 32'h00000000;
          16'h1ec1 : blkif.rom_rdata <= 32'h00000000;
          16'h1ec2 : blkif.rom_rdata <= 32'h00000000;
          16'h1ec3 : blkif.rom_rdata <= 32'h00000000;
          16'h1ec4 : blkif.rom_rdata <= 32'h00000000;
          16'h1ec5 : blkif.rom_rdata <= 32'h00000000;
          16'h1ec6 : blkif.rom_rdata <= 32'h00000000;
          16'h1ec7 : blkif.rom_rdata <= 32'h00000000;
          16'h1ec8 : blkif.rom_rdata <= 32'h00000000;
          16'h1ec9 : blkif.rom_rdata <= 32'h00000000;
          16'h1eca : blkif.rom_rdata <= 32'h00000000;
          16'h1ecb : blkif.rom_rdata <= 32'h00000000;
          16'h1ecc : blkif.rom_rdata <= 32'h00000000;
          16'h1ecd : blkif.rom_rdata <= 32'h00000000;
          16'h1ece : blkif.rom_rdata <= 32'h00000000;
          16'h1ecf : blkif.rom_rdata <= 32'h00000000;
          16'h1ed0 : blkif.rom_rdata <= 32'h00000000;
          16'h1ed1 : blkif.rom_rdata <= 32'h00000000;
          16'h1ed2 : blkif.rom_rdata <= 32'h00000000;
          16'h1ed3 : blkif.rom_rdata <= 32'h00000000;
          16'h1ed4 : blkif.rom_rdata <= 32'h00000000;
          16'h1ed5 : blkif.rom_rdata <= 32'h00000000;
          16'h1ed6 : blkif.rom_rdata <= 32'h00000000;
          16'h1ed7 : blkif.rom_rdata <= 32'h00000000;
          16'h1ed8 : blkif.rom_rdata <= 32'h00000000;
          16'h1ed9 : blkif.rom_rdata <= 32'h00000000;
          16'h1eda : blkif.rom_rdata <= 32'h00000000;
          16'h1edb : blkif.rom_rdata <= 32'h00000000;
          16'h1edc : blkif.rom_rdata <= 32'h00000000;
          16'h1edd : blkif.rom_rdata <= 32'h00000000;
          16'h1ede : blkif.rom_rdata <= 32'h00000000;
          16'h1edf : blkif.rom_rdata <= 32'h00000000;
          16'h1ee0 : blkif.rom_rdata <= 32'h00000000;
          16'h1ee1 : blkif.rom_rdata <= 32'h00000000;
          16'h1ee2 : blkif.rom_rdata <= 32'h00000000;
          16'h1ee3 : blkif.rom_rdata <= 32'h00000000;
          16'h1ee4 : blkif.rom_rdata <= 32'h00000000;
          16'h1ee5 : blkif.rom_rdata <= 32'h00000000;
          16'h1ee6 : blkif.rom_rdata <= 32'h00000000;
          16'h1ee7 : blkif.rom_rdata <= 32'h00000000;
          16'h1ee8 : blkif.rom_rdata <= 32'h00000000;
          16'h1ee9 : blkif.rom_rdata <= 32'h00000000;
          16'h1eea : blkif.rom_rdata <= 32'h00000000;
          16'h1eeb : blkif.rom_rdata <= 32'h00000000;
          16'h1eec : blkif.rom_rdata <= 32'h00000000;
          16'h1eed : blkif.rom_rdata <= 32'h00000000;
          16'h1eee : blkif.rom_rdata <= 32'h00000000;
          16'h1eef : blkif.rom_rdata <= 32'h00000000;
          16'h1ef0 : blkif.rom_rdata <= 32'h00000000;
          16'h1ef1 : blkif.rom_rdata <= 32'h00000000;
          16'h1ef2 : blkif.rom_rdata <= 32'h00000000;
          16'h1ef3 : blkif.rom_rdata <= 32'h00000000;
          16'h1ef4 : blkif.rom_rdata <= 32'h00000000;
          16'h1ef5 : blkif.rom_rdata <= 32'h00000000;
          16'h1ef6 : blkif.rom_rdata <= 32'h00000000;
          16'h1ef7 : blkif.rom_rdata <= 32'h00000000;
          16'h1ef8 : blkif.rom_rdata <= 32'h00000000;
          16'h1ef9 : blkif.rom_rdata <= 32'h00000000;
          16'h1efa : blkif.rom_rdata <= 32'h00000000;
          16'h1efb : blkif.rom_rdata <= 32'h00000000;
          16'h1efc : blkif.rom_rdata <= 32'h00000000;
          16'h1efd : blkif.rom_rdata <= 32'h00000000;
          16'h1efe : blkif.rom_rdata <= 32'h00000000;
          16'h1eff : blkif.rom_rdata <= 32'h00000000;
          16'h1f00 : blkif.rom_rdata <= 32'h00000000;
          16'h1f01 : blkif.rom_rdata <= 32'h00000000;
          16'h1f02 : blkif.rom_rdata <= 32'h00000000;
          16'h1f03 : blkif.rom_rdata <= 32'h00000000;
          16'h1f04 : blkif.rom_rdata <= 32'h00000000;
          16'h1f05 : blkif.rom_rdata <= 32'h00000000;
          16'h1f06 : blkif.rom_rdata <= 32'h00000000;
          16'h1f07 : blkif.rom_rdata <= 32'h00000000;
          16'h1f08 : blkif.rom_rdata <= 32'h00000000;
          16'h1f09 : blkif.rom_rdata <= 32'h00000000;
          16'h1f0a : blkif.rom_rdata <= 32'h00000000;
          16'h1f0b : blkif.rom_rdata <= 32'h00000000;
          16'h1f0c : blkif.rom_rdata <= 32'h00000000;
          16'h1f0d : blkif.rom_rdata <= 32'h00000000;
          16'h1f0e : blkif.rom_rdata <= 32'h00000000;
          16'h1f0f : blkif.rom_rdata <= 32'h00000000;
          16'h1f10 : blkif.rom_rdata <= 32'h00000000;
          16'h1f11 : blkif.rom_rdata <= 32'h00000000;
          16'h1f12 : blkif.rom_rdata <= 32'h00000000;
          16'h1f13 : blkif.rom_rdata <= 32'h00000000;
          16'h1f14 : blkif.rom_rdata <= 32'h00000000;
          16'h1f15 : blkif.rom_rdata <= 32'h00000000;
          16'h1f16 : blkif.rom_rdata <= 32'h00000000;
          16'h1f17 : blkif.rom_rdata <= 32'h00000000;
          16'h1f18 : blkif.rom_rdata <= 32'h00000000;
          16'h1f19 : blkif.rom_rdata <= 32'h00000000;
          16'h1f1a : blkif.rom_rdata <= 32'h00000000;
          16'h1f1b : blkif.rom_rdata <= 32'h00000000;
          16'h1f1c : blkif.rom_rdata <= 32'h00000000;
          16'h1f1d : blkif.rom_rdata <= 32'h00000000;
          16'h1f1e : blkif.rom_rdata <= 32'h00000000;
          16'h1f1f : blkif.rom_rdata <= 32'h00000000;
          16'h1f20 : blkif.rom_rdata <= 32'h00000000;
          16'h1f21 : blkif.rom_rdata <= 32'h00000000;
          16'h1f22 : blkif.rom_rdata <= 32'h00000000;
          16'h1f23 : blkif.rom_rdata <= 32'h00000000;
          16'h1f24 : blkif.rom_rdata <= 32'h00000000;
          16'h1f25 : blkif.rom_rdata <= 32'h00000000;
          16'h1f26 : blkif.rom_rdata <= 32'h00000000;
          16'h1f27 : blkif.rom_rdata <= 32'h00000000;
          16'h1f28 : blkif.rom_rdata <= 32'h00000000;
          16'h1f29 : blkif.rom_rdata <= 32'h00000000;
          16'h1f2a : blkif.rom_rdata <= 32'h00000000;
          16'h1f2b : blkif.rom_rdata <= 32'h00000000;
          16'h1f2c : blkif.rom_rdata <= 32'h00000000;
          16'h1f2d : blkif.rom_rdata <= 32'h00000000;
          16'h1f2e : blkif.rom_rdata <= 32'h00000000;
          16'h1f2f : blkif.rom_rdata <= 32'h00000000;
          16'h1f30 : blkif.rom_rdata <= 32'h00000000;
          16'h1f31 : blkif.rom_rdata <= 32'h00000000;
          16'h1f32 : blkif.rom_rdata <= 32'h00000000;
          16'h1f33 : blkif.rom_rdata <= 32'h00000000;
          16'h1f34 : blkif.rom_rdata <= 32'h00000000;
          16'h1f35 : blkif.rom_rdata <= 32'h00000000;
          16'h1f36 : blkif.rom_rdata <= 32'h00000000;
          16'h1f37 : blkif.rom_rdata <= 32'h00000000;
          16'h1f38 : blkif.rom_rdata <= 32'h00000000;
          16'h1f39 : blkif.rom_rdata <= 32'h00000000;
          16'h1f3a : blkif.rom_rdata <= 32'h00000000;
          16'h1f3b : blkif.rom_rdata <= 32'h00000000;
          16'h1f3c : blkif.rom_rdata <= 32'h00000000;
          16'h1f3d : blkif.rom_rdata <= 32'h00000000;
          16'h1f3e : blkif.rom_rdata <= 32'h00000000;
          16'h1f3f : blkif.rom_rdata <= 32'h00000000;
          16'h1f40 : blkif.rom_rdata <= 32'h00000000;
          16'h1f41 : blkif.rom_rdata <= 32'h00000000;
          16'h1f42 : blkif.rom_rdata <= 32'h00000000;
          16'h1f43 : blkif.rom_rdata <= 32'h00000000;
          16'h1f44 : blkif.rom_rdata <= 32'h00000000;
          16'h1f45 : blkif.rom_rdata <= 32'h00000000;
          16'h1f46 : blkif.rom_rdata <= 32'h00000000;
          16'h1f47 : blkif.rom_rdata <= 32'h00000000;
          16'h1f48 : blkif.rom_rdata <= 32'h00000000;
          16'h1f49 : blkif.rom_rdata <= 32'h00000000;
          16'h1f4a : blkif.rom_rdata <= 32'h00000000;
          16'h1f4b : blkif.rom_rdata <= 32'h00000000;
          16'h1f4c : blkif.rom_rdata <= 32'h00000000;
          16'h1f4d : blkif.rom_rdata <= 32'h00000000;
          16'h1f4e : blkif.rom_rdata <= 32'h00000000;
          16'h1f4f : blkif.rom_rdata <= 32'h00000000;
          16'h1f50 : blkif.rom_rdata <= 32'h00000000;
          16'h1f51 : blkif.rom_rdata <= 32'h00000000;
          16'h1f52 : blkif.rom_rdata <= 32'h00000000;
          16'h1f53 : blkif.rom_rdata <= 32'h00000000;
          16'h1f54 : blkif.rom_rdata <= 32'h00000000;
          16'h1f55 : blkif.rom_rdata <= 32'h00000000;
          16'h1f56 : blkif.rom_rdata <= 32'h00000000;
          16'h1f57 : blkif.rom_rdata <= 32'h00000000;
          16'h1f58 : blkif.rom_rdata <= 32'h00000000;
          16'h1f59 : blkif.rom_rdata <= 32'h00000000;
          16'h1f5a : blkif.rom_rdata <= 32'h00000000;
          16'h1f5b : blkif.rom_rdata <= 32'h00000000;
          16'h1f5c : blkif.rom_rdata <= 32'h00000000;
          16'h1f5d : blkif.rom_rdata <= 32'h00000000;
          16'h1f5e : blkif.rom_rdata <= 32'h00000000;
          16'h1f5f : blkif.rom_rdata <= 32'h00000000;
          16'h1f60 : blkif.rom_rdata <= 32'h00000000;
          16'h1f61 : blkif.rom_rdata <= 32'h00000000;
          16'h1f62 : blkif.rom_rdata <= 32'h00000000;
          16'h1f63 : blkif.rom_rdata <= 32'h00000000;
          16'h1f64 : blkif.rom_rdata <= 32'h00000000;
          16'h1f65 : blkif.rom_rdata <= 32'h00000000;
          16'h1f66 : blkif.rom_rdata <= 32'h00000000;
          16'h1f67 : blkif.rom_rdata <= 32'h00000000;
          16'h1f68 : blkif.rom_rdata <= 32'h00000000;
          16'h1f69 : blkif.rom_rdata <= 32'h00000000;
          16'h1f6a : blkif.rom_rdata <= 32'h00000000;
          16'h1f6b : blkif.rom_rdata <= 32'h00000000;
          16'h1f6c : blkif.rom_rdata <= 32'h00000000;
          16'h1f6d : blkif.rom_rdata <= 32'h00000000;
          16'h1f6e : blkif.rom_rdata <= 32'h00000000;
          16'h1f6f : blkif.rom_rdata <= 32'h00000000;
          16'h1f70 : blkif.rom_rdata <= 32'h00000000;
          16'h1f71 : blkif.rom_rdata <= 32'h00000000;
          16'h1f72 : blkif.rom_rdata <= 32'h00000000;
          16'h1f73 : blkif.rom_rdata <= 32'h00000000;
          16'h1f74 : blkif.rom_rdata <= 32'h00000000;
          16'h1f75 : blkif.rom_rdata <= 32'h00000000;
          16'h1f76 : blkif.rom_rdata <= 32'h00000000;
          16'h1f77 : blkif.rom_rdata <= 32'h00000000;
          16'h1f78 : blkif.rom_rdata <= 32'h00000000;
          16'h1f79 : blkif.rom_rdata <= 32'h00000000;
          16'h1f7a : blkif.rom_rdata <= 32'h00000000;
          16'h1f7b : blkif.rom_rdata <= 32'h00000000;
          16'h1f7c : blkif.rom_rdata <= 32'h00000000;
          16'h1f7d : blkif.rom_rdata <= 32'h00000000;
          16'h1f7e : blkif.rom_rdata <= 32'h00000000;
          16'h1f7f : blkif.rom_rdata <= 32'h00000000;
          16'h1f80 : blkif.rom_rdata <= 32'h00000000;
          16'h1f81 : blkif.rom_rdata <= 32'h00000000;
          16'h1f82 : blkif.rom_rdata <= 32'h00000000;
          16'h1f83 : blkif.rom_rdata <= 32'h00000000;
          16'h1f84 : blkif.rom_rdata <= 32'h00000000;
          16'h1f85 : blkif.rom_rdata <= 32'h00000000;
          16'h1f86 : blkif.rom_rdata <= 32'h00000000;
          16'h1f87 : blkif.rom_rdata <= 32'h00000000;
          16'h1f88 : blkif.rom_rdata <= 32'h00000000;
          16'h1f89 : blkif.rom_rdata <= 32'h00000000;
          16'h1f8a : blkif.rom_rdata <= 32'h00000000;
          16'h1f8b : blkif.rom_rdata <= 32'h00000000;
          16'h1f8c : blkif.rom_rdata <= 32'h00000000;
          16'h1f8d : blkif.rom_rdata <= 32'h00000000;
          16'h1f8e : blkif.rom_rdata <= 32'h00000000;
          16'h1f8f : blkif.rom_rdata <= 32'h00000000;
          16'h1f90 : blkif.rom_rdata <= 32'h00000000;
          16'h1f91 : blkif.rom_rdata <= 32'h00000000;
          16'h1f92 : blkif.rom_rdata <= 32'h00000000;
          16'h1f93 : blkif.rom_rdata <= 32'h00000000;
          16'h1f94 : blkif.rom_rdata <= 32'h00000000;
          16'h1f95 : blkif.rom_rdata <= 32'h00000000;
          16'h1f96 : blkif.rom_rdata <= 32'h00000000;
          16'h1f97 : blkif.rom_rdata <= 32'h00000000;
          16'h1f98 : blkif.rom_rdata <= 32'h00000000;
          16'h1f99 : blkif.rom_rdata <= 32'h00000000;
          16'h1f9a : blkif.rom_rdata <= 32'h00000000;
          16'h1f9b : blkif.rom_rdata <= 32'h00000000;
          16'h1f9c : blkif.rom_rdata <= 32'h00000000;
          16'h1f9d : blkif.rom_rdata <= 32'h00000000;
          16'h1f9e : blkif.rom_rdata <= 32'h00000000;
          16'h1f9f : blkif.rom_rdata <= 32'h00000000;
          16'h1fa0 : blkif.rom_rdata <= 32'h00000000;
          16'h1fa1 : blkif.rom_rdata <= 32'h00000000;
          16'h1fa2 : blkif.rom_rdata <= 32'h00000000;
          16'h1fa3 : blkif.rom_rdata <= 32'h00000000;
          16'h1fa4 : blkif.rom_rdata <= 32'h00000000;
          16'h1fa5 : blkif.rom_rdata <= 32'h00000000;
          16'h1fa6 : blkif.rom_rdata <= 32'h00000000;
          16'h1fa7 : blkif.rom_rdata <= 32'h00000000;
          16'h1fa8 : blkif.rom_rdata <= 32'h00000000;
          16'h1fa9 : blkif.rom_rdata <= 32'h00000000;
          16'h1faa : blkif.rom_rdata <= 32'h00000000;
          16'h1fab : blkif.rom_rdata <= 32'h00000000;
          16'h1fac : blkif.rom_rdata <= 32'h00000000;
          16'h1fad : blkif.rom_rdata <= 32'h00000000;
          16'h1fae : blkif.rom_rdata <= 32'h00000000;
          16'h1faf : blkif.rom_rdata <= 32'h00000000;
          16'h1fb0 : blkif.rom_rdata <= 32'h00000000;
          16'h1fb1 : blkif.rom_rdata <= 32'h00000000;
          16'h1fb2 : blkif.rom_rdata <= 32'h00000000;
          16'h1fb3 : blkif.rom_rdata <= 32'h00000000;
          16'h1fb4 : blkif.rom_rdata <= 32'h00000000;
          16'h1fb5 : blkif.rom_rdata <= 32'h00000000;
          16'h1fb6 : blkif.rom_rdata <= 32'h00000000;
          16'h1fb7 : blkif.rom_rdata <= 32'h00000000;
          16'h1fb8 : blkif.rom_rdata <= 32'h00000000;
          16'h1fb9 : blkif.rom_rdata <= 32'h00000000;
          16'h1fba : blkif.rom_rdata <= 32'h00000000;
          16'h1fbb : blkif.rom_rdata <= 32'h00000000;
          16'h1fbc : blkif.rom_rdata <= 32'h00000000;
          16'h1fbd : blkif.rom_rdata <= 32'h00000000;
          16'h1fbe : blkif.rom_rdata <= 32'h00000000;
          16'h1fbf : blkif.rom_rdata <= 32'h00000000;
          16'h1fc0 : blkif.rom_rdata <= 32'h00000000;
          16'h1fc1 : blkif.rom_rdata <= 32'h00000000;
          16'h1fc2 : blkif.rom_rdata <= 32'h00000000;
          16'h1fc3 : blkif.rom_rdata <= 32'h00000000;
          16'h1fc4 : blkif.rom_rdata <= 32'h00000000;
          16'h1fc5 : blkif.rom_rdata <= 32'h00000000;
          16'h1fc6 : blkif.rom_rdata <= 32'h00000000;
          16'h1fc7 : blkif.rom_rdata <= 32'h00000000;
          16'h1fc8 : blkif.rom_rdata <= 32'h00000000;
          16'h1fc9 : blkif.rom_rdata <= 32'h00000000;
          16'h1fca : blkif.rom_rdata <= 32'h00000000;
          16'h1fcb : blkif.rom_rdata <= 32'h00000000;
          16'h1fcc : blkif.rom_rdata <= 32'h00000000;
          16'h1fcd : blkif.rom_rdata <= 32'h00000000;
          16'h1fce : blkif.rom_rdata <= 32'h00000000;
          16'h1fcf : blkif.rom_rdata <= 32'h00000000;
          16'h1fd0 : blkif.rom_rdata <= 32'h00000000;
          16'h1fd1 : blkif.rom_rdata <= 32'h00000000;
          16'h1fd2 : blkif.rom_rdata <= 32'h00000000;
          16'h1fd3 : blkif.rom_rdata <= 32'h00000000;
          16'h1fd4 : blkif.rom_rdata <= 32'h00000000;
          16'h1fd5 : blkif.rom_rdata <= 32'h00000000;
          16'h1fd6 : blkif.rom_rdata <= 32'h00000000;
          16'h1fd7 : blkif.rom_rdata <= 32'h00000000;
          16'h1fd8 : blkif.rom_rdata <= 32'h00000000;
          16'h1fd9 : blkif.rom_rdata <= 32'h00000000;
          16'h1fda : blkif.rom_rdata <= 32'h00000000;
          16'h1fdb : blkif.rom_rdata <= 32'h00000000;
          16'h1fdc : blkif.rom_rdata <= 32'h00000000;
          16'h1fdd : blkif.rom_rdata <= 32'h00000000;
          16'h1fde : blkif.rom_rdata <= 32'h00000000;
          16'h1fdf : blkif.rom_rdata <= 32'h00000000;
          16'h1fe0 : blkif.rom_rdata <= 32'h00000000;
          16'h1fe1 : blkif.rom_rdata <= 32'h00000000;
          16'h1fe2 : blkif.rom_rdata <= 32'h00000000;
          16'h1fe3 : blkif.rom_rdata <= 32'h00000000;
          16'h1fe4 : blkif.rom_rdata <= 32'h00000000;
          16'h1fe5 : blkif.rom_rdata <= 32'h00000000;
          16'h1fe6 : blkif.rom_rdata <= 32'h00000000;
          16'h1fe7 : blkif.rom_rdata <= 32'h00000000;
          16'h1fe8 : blkif.rom_rdata <= 32'h00000000;
          16'h1fe9 : blkif.rom_rdata <= 32'h00000000;
          16'h1fea : blkif.rom_rdata <= 32'h00000000;
          16'h1feb : blkif.rom_rdata <= 32'h00000000;
          16'h1fec : blkif.rom_rdata <= 32'h00000000;
          16'h1fed : blkif.rom_rdata <= 32'h00000000;
          16'h1fee : blkif.rom_rdata <= 32'h00000000;
          16'h1fef : blkif.rom_rdata <= 32'h00000000;
          16'h1ff0 : blkif.rom_rdata <= 32'h00000000;
          16'h1ff1 : blkif.rom_rdata <= 32'h00000000;
          16'h1ff2 : blkif.rom_rdata <= 32'h00000000;
          16'h1ff3 : blkif.rom_rdata <= 32'h00000000;
          16'h1ff4 : blkif.rom_rdata <= 32'h00000000;
          16'h1ff5 : blkif.rom_rdata <= 32'h00000000;
          16'h1ff6 : blkif.rom_rdata <= 32'h00000000;
          16'h1ff7 : blkif.rom_rdata <= 32'h00000000;
          16'h1ff8 : blkif.rom_rdata <= 32'h00000000;
          16'h1ff9 : blkif.rom_rdata <= 32'h00000000;
          16'h1ffa : blkif.rom_rdata <= 32'h00000000;
          16'h1ffb : blkif.rom_rdata <= 32'h00000000;
          16'h1ffc : blkif.rom_rdata <= 32'h00000000;
          16'h1ffd : blkif.rom_rdata <= 32'h00000000;
          16'h1ffe : blkif.rom_rdata <= 32'h00000000;
          16'h1fff : blkif.rom_rdata <= 32'h00000000;
          default : blkif.rom_rdata <= 32'hDEADBEEF;
        endcase
end
endmodule

