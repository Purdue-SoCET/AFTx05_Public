module Memory_RAO
#(parameter integer ADDRBITSIZE = 16,parameter integer DATABITSIZE = 32,parameter integer TOPROM = 16)
(input wire clk,input wire n_rst,input wire [DATABITSIZE - 1:0] w_data,input wire [ADDRBITSIZE - 1:0] addr,input wire w_en,output reg [DATABITSIZE - 1:0] data);
reg [DATABITSIZE - 1:0] TOPRAMdata;		//RAM Data
reg [DATABITSIZE - 1:0] BOTTOMRAMdata;	//RAM Data
logic [ADDRBITSIZE - 1:0] reg_addr;
logic topw_en;
 logic unsigned [ADDRBITSIZE - 1:0] addr_top;
always_ff @(posedge clk) begin reg_addr <= addr; end
	SOC_RAM #(.ADDRBIT(ADDRBITSIZE),.DATABIT(DATABITSIZE),.BOTTOMADDR(0),.TOPADDR(128)) TOPRAM(.clk(clk),.n_rst(n_rst),.w_data(w_data),.addr(addr_top),.w_en(topw_en),.r_data(TOPRAMdata));
	SOC_RAM #(.ADDRBIT(ADDRBITSIZE),.DATABIT(DATABITSIZE),.BOTTOMADDR(0),.TOPADDR(58)) BOTTOMRAM(.clk(clk),.n_rst(n_rst),.w_data(w_data),.addr(addr),.w_en(w_en),.r_data(BOTTOMRAMdata));
assign addr_top = addr - 16'h2db3;
always_comb begin if((reg_addr < (16'h3b))) begin data <= BOTTOMRAMdata; end
else if (reg_addr < (16'h2db3)) begin case (reg_addr)
	16'h3b : data <= 32'h00020000;
	16'h3f : data <= 32'h03000000;
	16'h40 : data <= 32'h178f0000;
	16'h41 : data <= 32'h130f4f97;
	16'h42 : data <= 32'hf32f1034;
	16'h43 : data <= 32'h630cff07;
	16'h44 : data <= 32'h170f0000;
	16'h45 : data <= 32'h130f0fef;
	16'h46 : data <= 32'h63180f02;
	16'h47 : data <= 32'h170f0000;
	16'h48 : data <= 32'h130f4fee;
	16'h49 : data <= 32'h63040f00;
	16'h4a : data <= 32'h6ff09fed;
	16'h4b : data <= 32'h6f004005;
	16'h4c : data <= 32'h13000000;
	16'h4d : data <= 32'h13000000;
	16'h4e : data <= 32'h13000000;
	16'h4f : data <= 32'h13000000;
	16'h50 : data <= 32'h732f2034;
	16'h51 : data <= 32'he35e0ffa;
	16'h52 : data <= 32'h73005030;
	16'h53 : data <= 32'h13000000;
	16'h54 : data <= 32'h13000000;
	16'h55 : data <= 32'h13000000;
	16'h56 : data <= 32'h13000000;
	16'h57 : data <= 32'h13000000;
	16'h58 : data <= 32'h13000000;
	16'h59 : data <= 32'h13000000;
	16'h5a : data <= 32'h13000000;
	16'h5b : data <= 32'h13000000;
	16'h5c : data <= 32'h13000000;
	16'h5d : data <= 32'h13000000;
	16'h5e : data <= 32'h13000000;
	16'h5f : data <= 32'h13000000;
	16'h60 : data <= 32'h136e9e53;
	16'h61 : data <= 32'h73100e78;
	16'h62 : data <= 32'h6ff0dfff;
	16'h63 : data <= 32'h13000000;
	16'h64 : data <= 32'h13000000;
	16'h65 : data <= 32'h13000000;
	16'h66 : data <= 32'h13000000;
	16'h67 : data <= 32'h13000000;
	16'h68 : data <= 32'h13000000;
	16'h69 : data <= 32'h13000000;
	16'h6a : data <= 32'h13000000;
	16'h6b : data <= 32'h13000000;
	16'h6c : data <= 32'h13000000;
	16'h6d : data <= 32'h13000000;
	16'h6e : data <= 32'h13000000;
	16'h6f : data <= 32'h13000000;
	16'h70 : data <= 32'h178f0000;
	16'h71 : data <= 32'h130f4f8b;
	16'h72 : data <= 32'hf32f1034;
	16'h73 : data <= 32'he30cfffb;
	16'h74 : data <= 32'h170f0000;
	16'h75 : data <= 32'h130f0fe3;
	16'h76 : data <= 32'h63040f00;
	16'h77 : data <= 32'h6ff05fe2;
	16'h78 : data <= 32'h6ff01ffa;
	16'h79 : data <= 32'h13000000;
	16'h7a : data <= 32'h13000000;
	16'h7b : data <= 32'h13000000;
	16'h7c : data <= 32'h13000000;
	16'h7d : data <= 32'h13000000;
	16'h7e : data <= 32'h13000000;
	16'h7f : data <= 32'h13000000;
	16'h80 : data <= 32'h732500f1;
	16'h81 : data <= 32'h63100500;
	16'h82 : data <= 32'h732500f0;
	16'h83 : data <= 32'h63580500;
	16'h84 : data <= 32'h0f00f00f;
	16'h85 : data <= 32'h130e1000;
	16'h86 : data <= 32'h6f70d005;
	16'h87 : data <= 32'h97020000;
	16'h88 : data <= 32'h938242de;
	16'h89 : data <= 32'h63840200;
	16'h8a : data <= 32'h73901210;
	16'h8b : data <= 32'h9302801f;
	16'h8c : data <= 32'h73b00230;
	16'h8d : data <= 32'h97020000;
	16'h8e : data <= 32'h93824201;
	16'h8f : data <= 32'h73901234;
	16'h90 : data <= 32'h732500f1;
	16'h91 : data <= 32'h73000010;
	16'h92 : data <= 32'hb7000080;
	16'h93 : data <= 32'h93804000;
	16'h94 : data <= 32'h37010100;
	16'h95 : data <= 32'h1301f1ff;
	16'h96 : data <= 32'h23a02000;
	16'h97 : data <= 32'h37c10000;
	16'h98 : data <= 32'h1301f1ee;
	16'h99 : data <= 32'hb7000080;
	16'h9a : data <= 32'h93808000;
	16'h9b : data <= 32'h23a02000;
	16'h9c : data <= 32'h93000000;
	16'h9d : data <= 32'h13010000;
	16'h9e : data <= 32'hb3812000;
	16'h9f : data <= 32'h930e0000;
	16'ha0 : data <= 32'h130e2000;
	16'ha1 : data <= 32'h6384d101;
	16'ha2 : data <= 32'h6f70c07c;
	16'ha3 : data <= 32'h93001000;
	16'ha4 : data <= 32'h13011000;
	16'ha5 : data <= 32'hb3812000;
	16'ha6 : data <= 32'h930e2000;
	16'ha7 : data <= 32'h130e3000;
	16'ha8 : data <= 32'h6384d101;
	16'ha9 : data <= 32'h6f70007b;
	16'haa : data <= 32'h93003000;
	16'hab : data <= 32'h13017000;
	16'hac : data <= 32'hb3812000;
	16'had : data <= 32'h930ea000;
	16'hae : data <= 32'h130e4000;
	16'haf : data <= 32'h6384d101;
	16'hb0 : data <= 32'h6f704079;
	16'hb1 : data <= 32'h93000000;
	16'hb2 : data <= 32'h3781ffff;
	16'hb3 : data <= 32'hb3812000;
	16'hb4 : data <= 32'hb78effff;
	16'hb5 : data <= 32'h130e5000;
	16'hb6 : data <= 32'h6384d101;
	16'hb7 : data <= 32'h6f708077;
	16'hb8 : data <= 32'hb7000080;
	16'hb9 : data <= 32'h13010000;
	16'hba : data <= 32'hb3812000;
	16'hbb : data <= 32'hb70e0080;
	16'hbc : data <= 32'h130e6000;
	16'hbd : data <= 32'h6384d101;
	16'hbe : data <= 32'h6f70c075;
	16'hbf : data <= 32'hb7000080;
	16'hc0 : data <= 32'h3781ffff;
	16'hc1 : data <= 32'hb3812000;
	16'hc2 : data <= 32'hb78eff7f;
	16'hc3 : data <= 32'h130e7000;
	16'hc4 : data <= 32'h6384d101;
	16'hc5 : data <= 32'h6f700074;
	16'hc6 : data <= 32'h93000000;
	16'hc7 : data <= 32'h37810000;
	16'hc8 : data <= 32'h1301f1ff;
	16'hc9 : data <= 32'hb3812000;
	16'hca : data <= 32'hb78e0000;
	16'hcb : data <= 32'h938efeff;
	16'hcc : data <= 32'h130e8000;
	16'hcd : data <= 32'h6384d101;
	16'hce : data <= 32'h6f70c071;
	16'hcf : data <= 32'hb7000080;
	16'hd0 : data <= 32'h9380f0ff;
	16'hd1 : data <= 32'h13010000;
	16'hd2 : data <= 32'hb3812000;
	16'hd3 : data <= 32'hb70e0080;
	16'hd4 : data <= 32'h938efeff;
	16'hd5 : data <= 32'h130e9000;
	16'hd6 : data <= 32'h6384d101;
	16'hd7 : data <= 32'h6f70806f;
	16'hd8 : data <= 32'hb7000080;
	16'hd9 : data <= 32'h9380f0ff;
	16'hda : data <= 32'h37810000;
	16'hdb : data <= 32'h1301f1ff;
	16'hdc : data <= 32'hb3812000;
	16'hdd : data <= 32'hb78e0080;
	16'hde : data <= 32'h938eeeff;
	16'hdf : data <= 32'h130ea000;
	16'he0 : data <= 32'h6384d101;
	16'he1 : data <= 32'h6f70006d;
	16'he2 : data <= 32'hb7000080;
	16'he3 : data <= 32'h37810000;
	16'he4 : data <= 32'h1301f1ff;
	16'he5 : data <= 32'hb3812000;
	16'he6 : data <= 32'hb78e0080;
	16'he7 : data <= 32'h938efeff;
	16'he8 : data <= 32'h130eb000;
	16'he9 : data <= 32'h6384d101;
	16'hea : data <= 32'h6f70c06a;
	16'heb : data <= 32'hb7000080;
	16'hec : data <= 32'h9380f0ff;
	16'hed : data <= 32'h3781ffff;
	16'hee : data <= 32'hb3812000;
	16'hef : data <= 32'hb78eff7f;
	16'hf0 : data <= 32'h938efeff;
	16'hf1 : data <= 32'h130ec000;
	16'hf2 : data <= 32'h6384d101;
	16'hf3 : data <= 32'h6f708068;
	16'hf4 : data <= 32'h93000000;
	16'hf5 : data <= 32'h1301f0ff;
	16'hf6 : data <= 32'hb3812000;
	16'hf7 : data <= 32'h930ef0ff;
	16'hf8 : data <= 32'h130ed000;
	16'hf9 : data <= 32'h6384d101;
	16'hfa : data <= 32'h6f70c066;
	16'hfb : data <= 32'h9300f0ff;
	16'hfc : data <= 32'h13011000;
	16'hfd : data <= 32'hb3812000;
	16'hfe : data <= 32'h930e0000;
	16'hff : data <= 32'h130ee000;
	16'h100 : data <= 32'h6384d101;
	16'h101 : data <= 32'h6f700065;
	16'h102 : data <= 32'h9300f0ff;
	16'h103 : data <= 32'h1301f0ff;
	16'h104 : data <= 32'hb3812000;
	16'h105 : data <= 32'h930ee0ff;
	16'h106 : data <= 32'h130ef000;
	16'h107 : data <= 32'h6384d101;
	16'h108 : data <= 32'h6f704063;
	16'h109 : data <= 32'h93001000;
	16'h10a : data <= 32'h37010080;
	16'h10b : data <= 32'h1301f1ff;
	16'h10c : data <= 32'hb3812000;
	16'h10d : data <= 32'hb70e0080;
	16'h10e : data <= 32'h130e0001;
	16'h10f : data <= 32'h6384d101;
	16'h110 : data <= 32'h6f704061;
	16'h111 : data <= 32'h9300d000;
	16'h112 : data <= 32'h1301b000;
	16'h113 : data <= 32'hb3802000;
	16'h114 : data <= 32'h930e8001;
	16'h115 : data <= 32'h130e1001;
	16'h116 : data <= 32'h6384d001;
	16'h117 : data <= 32'h6f70805f;
	16'h118 : data <= 32'h9300e000;
	16'h119 : data <= 32'h1301b000;
	16'h11a : data <= 32'h33812000;
	16'h11b : data <= 32'h930e9001;
	16'h11c : data <= 32'h130e2001;
	16'h11d : data <= 32'h6304d101;
	16'h11e : data <= 32'h6f70c05d;
	16'h11f : data <= 32'h9300d000;
	16'h120 : data <= 32'hb3801000;
	16'h121 : data <= 32'h930ea001;
	16'h122 : data <= 32'h130e3001;
	16'h123 : data <= 32'h6384d001;
	16'h124 : data <= 32'h6f70405c;
	16'h125 : data <= 32'h13020000;
	16'h126 : data <= 32'h9300d000;
	16'h127 : data <= 32'h1301b000;
	16'h128 : data <= 32'hb3812000;
	16'h129 : data <= 32'h13830100;
	16'h12a : data <= 32'h13021200;
	16'h12b : data <= 32'h93022000;
	16'h12c : data <= 32'he31452fe;
	16'h12d : data <= 32'h930e8001;
	16'h12e : data <= 32'h130e4001;
	16'h12f : data <= 32'h6304d301;
	16'h130 : data <= 32'h6f704059;
	16'h131 : data <= 32'h13020000;
	16'h132 : data <= 32'h9300e000;
	16'h133 : data <= 32'h1301b000;
	16'h134 : data <= 32'hb3812000;
	16'h135 : data <= 32'h13000000;
	16'h136 : data <= 32'h13830100;
	16'h137 : data <= 32'h13021200;
	16'h138 : data <= 32'h93022000;
	16'h139 : data <= 32'he31252fe;
	16'h13a : data <= 32'h930e9001;
	16'h13b : data <= 32'h130e5001;
	16'h13c : data <= 32'h6304d301;
	16'h13d : data <= 32'h6f700056;
	16'h13e : data <= 32'h13020000;
	16'h13f : data <= 32'h9300f000;
	16'h140 : data <= 32'h1301b000;
	16'h141 : data <= 32'hb3812000;
	16'h142 : data <= 32'h13000000;
	16'h143 : data <= 32'h13000000;
	16'h144 : data <= 32'h13830100;
	16'h145 : data <= 32'h13021200;
	16'h146 : data <= 32'h93022000;
	16'h147 : data <= 32'he31052fe;
	16'h148 : data <= 32'h930ea001;
	16'h149 : data <= 32'h130e6001;
	16'h14a : data <= 32'h6304d301;
	16'h14b : data <= 32'h6f708052;
	16'h14c : data <= 32'h13020000;
	16'h14d : data <= 32'h9300d000;
	16'h14e : data <= 32'h1301b000;
	16'h14f : data <= 32'hb3812000;
	16'h150 : data <= 32'h13021200;
	16'h151 : data <= 32'h93022000;
	16'h152 : data <= 32'he31652fe;
	16'h153 : data <= 32'h930e8001;
	16'h154 : data <= 32'h130e7001;
	16'h155 : data <= 32'h6384d101;
	16'h156 : data <= 32'h6f70c04f;
	16'h157 : data <= 32'h13020000;
	16'h158 : data <= 32'h9300e000;
	16'h159 : data <= 32'h1301b000;
	16'h15a : data <= 32'h13000000;
	16'h15b : data <= 32'hb3812000;
	16'h15c : data <= 32'h13021200;
	16'h15d : data <= 32'h93022000;
	16'h15e : data <= 32'he31452fe;
	16'h15f : data <= 32'h930e9001;
	16'h160 : data <= 32'h130e8001;
	16'h161 : data <= 32'h6384d101;
	16'h162 : data <= 32'h6f70c04c;
	16'h163 : data <= 32'h13020000;
	16'h164 : data <= 32'h9300f000;
	16'h165 : data <= 32'h1301b000;
	16'h166 : data <= 32'h13000000;
	16'h167 : data <= 32'h13000000;
	16'h168 : data <= 32'hb3812000;
	16'h169 : data <= 32'h13021200;
	16'h16a : data <= 32'h93022000;
	16'h16b : data <= 32'he31252fe;
	16'h16c : data <= 32'h930ea001;
	16'h16d : data <= 32'h130e9001;
	16'h16e : data <= 32'h6384d101;
	16'h16f : data <= 32'h6f708049;
	16'h170 : data <= 32'h13020000;
	16'h171 : data <= 32'h9300d000;
	16'h172 : data <= 32'h13000000;
	16'h173 : data <= 32'h1301b000;
	16'h174 : data <= 32'hb3812000;
	16'h175 : data <= 32'h13021200;
	16'h176 : data <= 32'h93022000;
	16'h177 : data <= 32'he31452fe;
	16'h178 : data <= 32'h930e8001;
	16'h179 : data <= 32'h130ea001;
	16'h17a : data <= 32'h6384d101;
	16'h17b : data <= 32'h6f708046;
	16'h17c : data <= 32'h13020000;
	16'h17d : data <= 32'h9300e000;
	16'h17e : data <= 32'h13000000;
	16'h17f : data <= 32'h1301b000;
	16'h180 : data <= 32'h13000000;
	16'h181 : data <= 32'hb3812000;
	16'h182 : data <= 32'h13021200;
	16'h183 : data <= 32'h93022000;
	16'h184 : data <= 32'he31252fe;
	16'h185 : data <= 32'h930e9001;
	16'h186 : data <= 32'h130eb001;
	16'h187 : data <= 32'h6384d101;
	16'h188 : data <= 32'h6f704043;
	16'h189 : data <= 32'h13020000;
	16'h18a : data <= 32'h9300f000;
	16'h18b : data <= 32'h13000000;
	16'h18c : data <= 32'h13000000;
	16'h18d : data <= 32'h1301b000;
	16'h18e : data <= 32'hb3812000;
	16'h18f : data <= 32'h13021200;
	16'h190 : data <= 32'h93022000;
	16'h191 : data <= 32'he31252fe;
	16'h192 : data <= 32'h930ea001;
	16'h193 : data <= 32'h130ec001;
	16'h194 : data <= 32'h6384d101;
	16'h195 : data <= 32'h6f700040;
	16'h196 : data <= 32'h13020000;
	16'h197 : data <= 32'h1301b000;
	16'h198 : data <= 32'h9300d000;
	16'h199 : data <= 32'hb3812000;
	16'h19a : data <= 32'h13021200;
	16'h19b : data <= 32'h93022000;
	16'h19c : data <= 32'he31652fe;
	16'h19d : data <= 32'h930e8001;
	16'h19e : data <= 32'h130ed001;
	16'h19f : data <= 32'h6384d101;
	16'h1a0 : data <= 32'h6f70403d;
	16'h1a1 : data <= 32'h13020000;
	16'h1a2 : data <= 32'h1301b000;
	16'h1a3 : data <= 32'h9300e000;
	16'h1a4 : data <= 32'h13000000;
	16'h1a5 : data <= 32'hb3812000;
	16'h1a6 : data <= 32'h13021200;
	16'h1a7 : data <= 32'h93022000;
	16'h1a8 : data <= 32'he31452fe;
	16'h1a9 : data <= 32'h930e9001;
	16'h1aa : data <= 32'h130ee001;
	16'h1ab : data <= 32'h6384d101;
	16'h1ac : data <= 32'h6f70403a;
	16'h1ad : data <= 32'h13020000;
	16'h1ae : data <= 32'h1301b000;
	16'h1af : data <= 32'h9300f000;
	16'h1b0 : data <= 32'h13000000;
	16'h1b1 : data <= 32'h13000000;
	16'h1b2 : data <= 32'hb3812000;
	16'h1b3 : data <= 32'h13021200;
	16'h1b4 : data <= 32'h93022000;
	16'h1b5 : data <= 32'he31252fe;
	16'h1b6 : data <= 32'h930ea001;
	16'h1b7 : data <= 32'h130ef001;
	16'h1b8 : data <= 32'h6384d101;
	16'h1b9 : data <= 32'h6f700037;
	16'h1ba : data <= 32'h13020000;
	16'h1bb : data <= 32'h1301b000;
	16'h1bc : data <= 32'h13000000;
	16'h1bd : data <= 32'h9300d000;
	16'h1be : data <= 32'hb3812000;
	16'h1bf : data <= 32'h13021200;
	16'h1c0 : data <= 32'h93022000;
	16'h1c1 : data <= 32'he31452fe;
	16'h1c2 : data <= 32'h930e8001;
	16'h1c3 : data <= 32'h130e0002;
	16'h1c4 : data <= 32'h6384d101;
	16'h1c5 : data <= 32'h6f700034;
	16'h1c6 : data <= 32'h13020000;
	16'h1c7 : data <= 32'h1301b000;
	16'h1c8 : data <= 32'h13000000;
	16'h1c9 : data <= 32'h9300e000;
	16'h1ca : data <= 32'h13000000;
	16'h1cb : data <= 32'hb3812000;
	16'h1cc : data <= 32'h13021200;
	16'h1cd : data <= 32'h93022000;
	16'h1ce : data <= 32'he31252fe;
	16'h1cf : data <= 32'h930e9001;
	16'h1d0 : data <= 32'h130e1002;
	16'h1d1 : data <= 32'h6384d101;
	16'h1d2 : data <= 32'h6f70c030;
	16'h1d3 : data <= 32'h13020000;
	16'h1d4 : data <= 32'h1301b000;
	16'h1d5 : data <= 32'h13000000;
	16'h1d6 : data <= 32'h13000000;
	16'h1d7 : data <= 32'h9300f000;
	16'h1d8 : data <= 32'hb3812000;
	16'h1d9 : data <= 32'h13021200;
	16'h1da : data <= 32'h93022000;
	16'h1db : data <= 32'he31252fe;
	16'h1dc : data <= 32'h930ea001;
	16'h1dd : data <= 32'h130e2002;
	16'h1de : data <= 32'h6384d101;
	16'h1df : data <= 32'h6f70802d;
	16'h1e0 : data <= 32'h9300f000;
	16'h1e1 : data <= 32'h33011000;
	16'h1e2 : data <= 32'h930ef000;
	16'h1e3 : data <= 32'h130e3002;
	16'h1e4 : data <= 32'h6304d101;
	16'h1e5 : data <= 32'h6f70002c;
	16'h1e6 : data <= 32'h93000002;
	16'h1e7 : data <= 32'h33810000;
	16'h1e8 : data <= 32'h930e0002;
	16'h1e9 : data <= 32'h130e4002;
	16'h1ea : data <= 32'h6304d101;
	16'h1eb : data <= 32'h6f70802a;
	16'h1ec : data <= 32'hb3000000;
	16'h1ed : data <= 32'h930e0000;
	16'h1ee : data <= 32'h130e5002;
	16'h1ef : data <= 32'h6384d001;
	16'h1f0 : data <= 32'h6f704029;
	16'h1f1 : data <= 32'h93000001;
	16'h1f2 : data <= 32'h1301e001;
	16'h1f3 : data <= 32'h33802000;
	16'h1f4 : data <= 32'h930e0000;
	16'h1f5 : data <= 32'h130e6002;
	16'h1f6 : data <= 32'h6304d001;
	16'h1f7 : data <= 32'h6f708027;
	16'h1f8 : data <= 32'h93000000;
	16'h1f9 : data <= 32'h93810000;
	16'h1fa : data <= 32'h930e0000;
	16'h1fb : data <= 32'h130e7002;
	16'h1fc : data <= 32'h6384d101;
	16'h1fd : data <= 32'h6f700026;
	16'h1fe : data <= 32'h93001000;
	16'h1ff : data <= 32'h93811000;
	16'h200 : data <= 32'h930e2000;
	16'h201 : data <= 32'h130e8002;
	16'h202 : data <= 32'h6384d101;
	16'h203 : data <= 32'h6f708024;
	16'h204 : data <= 32'h93003000;
	16'h205 : data <= 32'h93817000;
	16'h206 : data <= 32'h930ea000;
	16'h207 : data <= 32'h130e9002;
	16'h208 : data <= 32'h6384d101;
	16'h209 : data <= 32'h6f700023;
	16'h20a : data <= 32'h93000000;
	16'h20b : data <= 32'h93810080;
	16'h20c : data <= 32'h930e0080;
	16'h20d : data <= 32'h130ea002;
	16'h20e : data <= 32'h6384d101;
	16'h20f : data <= 32'h6f708021;
	16'h210 : data <= 32'hb7000080;
	16'h211 : data <= 32'h93810000;
	16'h212 : data <= 32'hb70e0080;
	16'h213 : data <= 32'h130eb002;
	16'h214 : data <= 32'h6384d101;
	16'h215 : data <= 32'h6f700020;
	16'h216 : data <= 32'hb7000080;
	16'h217 : data <= 32'h93810080;
	16'h218 : data <= 32'hb70e0080;
	16'h219 : data <= 32'h938e0e80;
	16'h21a : data <= 32'h130ec002;
	16'h21b : data <= 32'h6384d101;
	16'h21c : data <= 32'h6f70401e;
	16'h21d : data <= 32'h93000000;
	16'h21e : data <= 32'h9381f07f;
	16'h21f : data <= 32'h930ef07f;
	16'h220 : data <= 32'h130ed002;
	16'h221 : data <= 32'h6384d101;
	16'h222 : data <= 32'h6f70c01c;
	16'h223 : data <= 32'hb7000080;
	16'h224 : data <= 32'h9380f0ff;
	16'h225 : data <= 32'h93810000;
	16'h226 : data <= 32'hb70e0080;
	16'h227 : data <= 32'h938efeff;
	16'h228 : data <= 32'h130ee002;
	16'h229 : data <= 32'h6384d101;
	16'h22a : data <= 32'h6f70c01a;
	16'h22b : data <= 32'hb7000080;
	16'h22c : data <= 32'h9380f0ff;
	16'h22d : data <= 32'h9381f07f;
	16'h22e : data <= 32'hb70e0080;
	16'h22f : data <= 32'h938eee7f;
	16'h230 : data <= 32'h130ef002;
	16'h231 : data <= 32'h6384d101;
	16'h232 : data <= 32'h6f70c018;
	16'h233 : data <= 32'hb7000080;
	16'h234 : data <= 32'h9381f07f;
	16'h235 : data <= 32'hb70e0080;
	16'h236 : data <= 32'h938efe7f;
	16'h237 : data <= 32'h130e0003;
	16'h238 : data <= 32'h6384d101;
	16'h239 : data <= 32'h6f700017;
	16'h23a : data <= 32'hb7000080;
	16'h23b : data <= 32'h9380f0ff;
	16'h23c : data <= 32'h93810080;
	16'h23d : data <= 32'hb7feff7f;
	16'h23e : data <= 32'h938efe7f;
	16'h23f : data <= 32'h130e1003;
	16'h240 : data <= 32'h6384d101;
	16'h241 : data <= 32'h6f700015;
	16'h242 : data <= 32'h93000000;
	16'h243 : data <= 32'h9381f0ff;
	16'h244 : data <= 32'h930ef0ff;
	16'h245 : data <= 32'h130e2003;
	16'h246 : data <= 32'h6384d101;
	16'h247 : data <= 32'h6f708013;
	16'h248 : data <= 32'h9300f0ff;
	16'h249 : data <= 32'h93811000;
	16'h24a : data <= 32'h930e0000;
	16'h24b : data <= 32'h130e3003;
	16'h24c : data <= 32'h6384d101;
	16'h24d : data <= 32'h6f700012;
	16'h24e : data <= 32'h9300f0ff;
	16'h24f : data <= 32'h9381f0ff;
	16'h250 : data <= 32'h930ee0ff;
	16'h251 : data <= 32'h130e4003;
	16'h252 : data <= 32'h6384d101;
	16'h253 : data <= 32'h6f708010;
	16'h254 : data <= 32'hb7000080;
	16'h255 : data <= 32'h9380f0ff;
	16'h256 : data <= 32'h93811000;
	16'h257 : data <= 32'hb70e0080;
	16'h258 : data <= 32'h130e5003;
	16'h259 : data <= 32'h6384d101;
	16'h25a : data <= 32'h6f70c00e;
	16'h25b : data <= 32'h9300d000;
	16'h25c : data <= 32'h9380b000;
	16'h25d : data <= 32'h930e8001;
	16'h25e : data <= 32'h130e6003;
	16'h25f : data <= 32'h6384d001;
	16'h260 : data <= 32'h6f70400d;
	16'h261 : data <= 32'h13020000;
	16'h262 : data <= 32'h9300d000;
	16'h263 : data <= 32'h9381b000;
	16'h264 : data <= 32'h13830100;
	16'h265 : data <= 32'h13021200;
	16'h266 : data <= 32'h93022000;
	16'h267 : data <= 32'he31652fe;
	16'h268 : data <= 32'h930e8001;
	16'h269 : data <= 32'h130e7003;
	16'h26a : data <= 32'h6304d301;
	16'h26b : data <= 32'h6f70800a;
	16'h26c : data <= 32'h13020000;
	16'h26d : data <= 32'h9300d000;
	16'h26e : data <= 32'h9381a000;
	16'h26f : data <= 32'h13000000;
	16'h270 : data <= 32'h13830100;
	16'h271 : data <= 32'h13021200;
	16'h272 : data <= 32'h93022000;
	16'h273 : data <= 32'he31452fe;
	16'h274 : data <= 32'h930e7001;
	16'h275 : data <= 32'h130e8003;
	16'h276 : data <= 32'h6304d301;
	16'h277 : data <= 32'h6f708007;
	16'h278 : data <= 32'h13020000;
	16'h279 : data <= 32'h9300d000;
	16'h27a : data <= 32'h93819000;
	16'h27b : data <= 32'h13000000;
	16'h27c : data <= 32'h13000000;
	16'h27d : data <= 32'h13830100;
	16'h27e : data <= 32'h13021200;
	16'h27f : data <= 32'h93022000;
	16'h280 : data <= 32'he31252fe;
	16'h281 : data <= 32'h930e6001;
	16'h282 : data <= 32'h130e9003;
	16'h283 : data <= 32'h6304d301;
	16'h284 : data <= 32'h6f704004;
	16'h285 : data <= 32'h13020000;
	16'h286 : data <= 32'h9300d000;
	16'h287 : data <= 32'h9381b000;
	16'h288 : data <= 32'h13021200;
	16'h289 : data <= 32'h93022000;
	16'h28a : data <= 32'he31852fe;
	16'h28b : data <= 32'h930e8001;
	16'h28c : data <= 32'h130ea003;
	16'h28d : data <= 32'h6384d101;
	16'h28e : data <= 32'h6f70c001;
	16'h28f : data <= 32'h13020000;
	16'h290 : data <= 32'h9300d000;
	16'h291 : data <= 32'h13000000;
	16'h292 : data <= 32'h9381a000;
	16'h293 : data <= 32'h13021200;
	16'h294 : data <= 32'h93022000;
	16'h295 : data <= 32'he31652fe;
	16'h296 : data <= 32'h930e7001;
	16'h297 : data <= 32'h130eb003;
	16'h298 : data <= 32'h6384d101;
	16'h299 : data <= 32'h6f60107f;
	16'h29a : data <= 32'h13020000;
	16'h29b : data <= 32'h9300d000;
	16'h29c : data <= 32'h13000000;
	16'h29d : data <= 32'h13000000;
	16'h29e : data <= 32'h93819000;
	16'h29f : data <= 32'h13021200;
	16'h2a0 : data <= 32'h93022000;
	16'h2a1 : data <= 32'he31452fe;
	16'h2a2 : data <= 32'h930e6001;
	16'h2a3 : data <= 32'h130ec003;
	16'h2a4 : data <= 32'h6384d101;
	16'h2a5 : data <= 32'h6f60107c;
	16'h2a6 : data <= 32'h93000002;
	16'h2a7 : data <= 32'h930e0002;
	16'h2a8 : data <= 32'h130ed003;
	16'h2a9 : data <= 32'h6384d001;
	16'h2aa : data <= 32'h6f60d07a;
	16'h2ab : data <= 32'h93001002;
	16'h2ac : data <= 32'h13802003;
	16'h2ad : data <= 32'h930e0000;
	16'h2ae : data <= 32'h130ee003;
	16'h2af : data <= 32'h6304d001;
	16'h2b0 : data <= 32'h6f605079;
	16'h2b1 : data <= 32'hb70001ff;
	16'h2b2 : data <= 32'h938000f0;
	16'h2b3 : data <= 32'h37110f0f;
	16'h2b4 : data <= 32'h1301f1f0;
	16'h2b5 : data <= 32'hb3f12000;
	16'h2b6 : data <= 32'hb71e000f;
	16'h2b7 : data <= 32'h938e0ef0;
	16'h2b8 : data <= 32'h130ef003;
	16'h2b9 : data <= 32'h6384d101;
	16'h2ba : data <= 32'h6f60d076;
	16'h2bb : data <= 32'hb710f00f;
	16'h2bc : data <= 32'h938000ff;
	16'h2bd : data <= 32'h37f1f0f0;
	16'h2be : data <= 32'h1301010f;
	16'h2bf : data <= 32'hb3f12000;
	16'h2c0 : data <= 32'hb70ef000;
	16'h2c1 : data <= 32'h938e0e0f;
	16'h2c2 : data <= 32'h130e0004;
	16'h2c3 : data <= 32'h6384d101;
	16'h2c4 : data <= 32'h6f605074;
	16'h2c5 : data <= 32'hb700ff00;
	16'h2c6 : data <= 32'h9380f00f;
	16'h2c7 : data <= 32'h37110f0f;
	16'h2c8 : data <= 32'h1301f1f0;
	16'h2c9 : data <= 32'hb3f12000;
	16'h2ca : data <= 32'hb70e0f00;
	16'h2cb : data <= 32'h938efe00;
	16'h2cc : data <= 32'h130e1004;
	16'h2cd : data <= 32'h6384d101;
	16'h2ce : data <= 32'h6f60d071;
	16'h2cf : data <= 32'hb7f00ff0;
	16'h2d0 : data <= 32'h9380f000;
	16'h2d1 : data <= 32'h37f1f0f0;
	16'h2d2 : data <= 32'h1301010f;
	16'h2d3 : data <= 32'hb3f12000;
	16'h2d4 : data <= 32'hb7fe00f0;
	16'h2d5 : data <= 32'h130e2004;
	16'h2d6 : data <= 32'h6384d101;
	16'h2d7 : data <= 32'h6f60906f;
	16'h2d8 : data <= 32'hb70001ff;
	16'h2d9 : data <= 32'h938000f0;
	16'h2da : data <= 32'h37110f0f;
	16'h2db : data <= 32'h1301f1f0;
	16'h2dc : data <= 32'hb3f02000;
	16'h2dd : data <= 32'hb71e000f;
	16'h2de : data <= 32'h938e0ef0;
	16'h2df : data <= 32'h130e3004;
	16'h2e0 : data <= 32'h6384d001;
	16'h2e1 : data <= 32'h6f60106d;
	16'h2e2 : data <= 32'hb710f00f;
	16'h2e3 : data <= 32'h938000ff;
	16'h2e4 : data <= 32'h37f1f0f0;
	16'h2e5 : data <= 32'h1301010f;
	16'h2e6 : data <= 32'h33f12000;
	16'h2e7 : data <= 32'hb70ef000;
	16'h2e8 : data <= 32'h938e0e0f;
	16'h2e9 : data <= 32'h130e4004;
	16'h2ea : data <= 32'h6304d101;
	16'h2eb : data <= 32'h6f60906a;
	16'h2ec : data <= 32'hb70001ff;
	16'h2ed : data <= 32'h938000f0;
	16'h2ee : data <= 32'hb3f01000;
	16'h2ef : data <= 32'hb70e01ff;
	16'h2f0 : data <= 32'h938e0ef0;
	16'h2f1 : data <= 32'h130e5004;
	16'h2f2 : data <= 32'h6384d001;
	16'h2f3 : data <= 32'h6f609068;
	16'h2f4 : data <= 32'h13020000;
	16'h2f5 : data <= 32'hb70001ff;
	16'h2f6 : data <= 32'h938000f0;
	16'h2f7 : data <= 32'h37110f0f;
	16'h2f8 : data <= 32'h1301f1f0;
	16'h2f9 : data <= 32'hb3f12000;
	16'h2fa : data <= 32'h13830100;
	16'h2fb : data <= 32'h13021200;
	16'h2fc : data <= 32'h93022000;
	16'h2fd : data <= 32'he31052fe;
	16'h2fe : data <= 32'hb71e000f;
	16'h2ff : data <= 32'h938e0ef0;
	16'h300 : data <= 32'h130e6004;
	16'h301 : data <= 32'h6304d301;
	16'h302 : data <= 32'h6f60d064;
	16'h303 : data <= 32'h13020000;
	16'h304 : data <= 32'hb710f00f;
	16'h305 : data <= 32'h938000ff;
	16'h306 : data <= 32'h37f1f0f0;
	16'h307 : data <= 32'h1301010f;
	16'h308 : data <= 32'hb3f12000;
	16'h309 : data <= 32'h13000000;
	16'h30a : data <= 32'h13830100;
	16'h30b : data <= 32'h13021200;
	16'h30c : data <= 32'h93022000;
	16'h30d : data <= 32'he31e52fc;
	16'h30e : data <= 32'hb70ef000;
	16'h30f : data <= 32'h938e0e0f;
	16'h310 : data <= 32'h130e7004;
	16'h311 : data <= 32'h6304d301;
	16'h312 : data <= 32'h6f60d060;
	16'h313 : data <= 32'h13020000;
	16'h314 : data <= 32'hb700ff00;
	16'h315 : data <= 32'h9380f00f;
	16'h316 : data <= 32'h37110f0f;
	16'h317 : data <= 32'h1301f1f0;
	16'h318 : data <= 32'hb3f12000;
	16'h319 : data <= 32'h13000000;
	16'h31a : data <= 32'h13000000;
	16'h31b : data <= 32'h13830100;
	16'h31c : data <= 32'h13021200;
	16'h31d : data <= 32'h93022000;
	16'h31e : data <= 32'he31c52fc;
	16'h31f : data <= 32'hb70e0f00;
	16'h320 : data <= 32'h938efe00;
	16'h321 : data <= 32'h130e8004;
	16'h322 : data <= 32'h6304d301;
	16'h323 : data <= 32'h6f60905c;
	16'h324 : data <= 32'h13020000;
	16'h325 : data <= 32'hb70001ff;
	16'h326 : data <= 32'h938000f0;
	16'h327 : data <= 32'h37110f0f;
	16'h328 : data <= 32'h1301f1f0;
	16'h329 : data <= 32'hb3f12000;
	16'h32a : data <= 32'h13021200;
	16'h32b : data <= 32'h93022000;
	16'h32c : data <= 32'he31252fe;
	16'h32d : data <= 32'hb71e000f;
	16'h32e : data <= 32'h938e0ef0;
	16'h32f : data <= 32'h130e9004;
	16'h330 : data <= 32'h6384d101;
	16'h331 : data <= 32'h6f601059;
	16'h332 : data <= 32'h13020000;
	16'h333 : data <= 32'hb710f00f;
	16'h334 : data <= 32'h938000ff;
	16'h335 : data <= 32'h37f1f0f0;
	16'h336 : data <= 32'h1301010f;
	16'h337 : data <= 32'h13000000;
	16'h338 : data <= 32'hb3f12000;
	16'h339 : data <= 32'h13021200;
	16'h33a : data <= 32'h93022000;
	16'h33b : data <= 32'he31052fe;
	16'h33c : data <= 32'hb70ef000;
	16'h33d : data <= 32'h938e0e0f;
	16'h33e : data <= 32'h130ea004;
	16'h33f : data <= 32'h6384d101;
	16'h340 : data <= 32'h6f605055;
	16'h341 : data <= 32'h13020000;
	16'h342 : data <= 32'hb700ff00;
	16'h343 : data <= 32'h9380f00f;
	16'h344 : data <= 32'h37110f0f;
	16'h345 : data <= 32'h1301f1f0;
	16'h346 : data <= 32'h13000000;
	16'h347 : data <= 32'h13000000;
	16'h348 : data <= 32'hb3f12000;
	16'h349 : data <= 32'h13021200;
	16'h34a : data <= 32'h93022000;
	16'h34b : data <= 32'he31e52fc;
	16'h34c : data <= 32'hb70e0f00;
	16'h34d : data <= 32'h938efe00;
	16'h34e : data <= 32'h130eb004;
	16'h34f : data <= 32'h6384d101;
	16'h350 : data <= 32'h6f605051;
	16'h351 : data <= 32'h13020000;
	16'h352 : data <= 32'hb70001ff;
	16'h353 : data <= 32'h938000f0;
	16'h354 : data <= 32'h13000000;
	16'h355 : data <= 32'h37110f0f;
	16'h356 : data <= 32'h1301f1f0;
	16'h357 : data <= 32'hb3f12000;
	16'h358 : data <= 32'h13021200;
	16'h359 : data <= 32'h93022000;
	16'h35a : data <= 32'he31052fe;
	16'h35b : data <= 32'hb71e000f;
	16'h35c : data <= 32'h938e0ef0;
	16'h35d : data <= 32'h130ec004;
	16'h35e : data <= 32'h6384d101;
	16'h35f : data <= 32'h6f60904d;
	16'h360 : data <= 32'h13020000;
	16'h361 : data <= 32'hb710f00f;
	16'h362 : data <= 32'h938000ff;
	16'h363 : data <= 32'h13000000;
	16'h364 : data <= 32'h37f1f0f0;
	16'h365 : data <= 32'h1301010f;
	16'h366 : data <= 32'h13000000;
	16'h367 : data <= 32'hb3f12000;
	16'h368 : data <= 32'h13021200;
	16'h369 : data <= 32'h93022000;
	16'h36a : data <= 32'he31e52fc;
	16'h36b : data <= 32'hb70ef000;
	16'h36c : data <= 32'h938e0e0f;
	16'h36d : data <= 32'h130ed004;
	16'h36e : data <= 32'h6384d101;
	16'h36f : data <= 32'h6f609049;
	16'h370 : data <= 32'h13020000;
	16'h371 : data <= 32'hb700ff00;
	16'h372 : data <= 32'h9380f00f;
	16'h373 : data <= 32'h13000000;
	16'h374 : data <= 32'h13000000;
	16'h375 : data <= 32'h37110f0f;
	16'h376 : data <= 32'h1301f1f0;
	16'h377 : data <= 32'hb3f12000;
	16'h378 : data <= 32'h13021200;
	16'h379 : data <= 32'h93022000;
	16'h37a : data <= 32'he31e52fc;
	16'h37b : data <= 32'hb70e0f00;
	16'h37c : data <= 32'h938efe00;
	16'h37d : data <= 32'h130ee004;
	16'h37e : data <= 32'h6384d101;
	16'h37f : data <= 32'h6f609045;
	16'h380 : data <= 32'h13020000;
	16'h381 : data <= 32'h37110f0f;
	16'h382 : data <= 32'h1301f1f0;
	16'h383 : data <= 32'hb70001ff;
	16'h384 : data <= 32'h938000f0;
	16'h385 : data <= 32'hb3f12000;
	16'h386 : data <= 32'h13021200;
	16'h387 : data <= 32'h93022000;
	16'h388 : data <= 32'he31252fe;
	16'h389 : data <= 32'hb71e000f;
	16'h38a : data <= 32'h938e0ef0;
	16'h38b : data <= 32'h130ef004;
	16'h38c : data <= 32'h6384d101;
	16'h38d : data <= 32'h6f601042;
	16'h38e : data <= 32'h13020000;
	16'h38f : data <= 32'h37f1f0f0;
	16'h390 : data <= 32'h1301010f;
	16'h391 : data <= 32'hb710f00f;
	16'h392 : data <= 32'h938000ff;
	16'h393 : data <= 32'h13000000;
	16'h394 : data <= 32'hb3f12000;
	16'h395 : data <= 32'h13021200;
	16'h396 : data <= 32'h93022000;
	16'h397 : data <= 32'he31052fe;
	16'h398 : data <= 32'hb70ef000;
	16'h399 : data <= 32'h938e0e0f;
	16'h39a : data <= 32'h130e0005;
	16'h39b : data <= 32'h6384d101;
	16'h39c : data <= 32'h6f60503e;
	16'h39d : data <= 32'h13020000;
	16'h39e : data <= 32'h37110f0f;
	16'h39f : data <= 32'h1301f1f0;
	16'h3a0 : data <= 32'hb700ff00;
	16'h3a1 : data <= 32'h9380f00f;
	16'h3a2 : data <= 32'h13000000;
	16'h3a3 : data <= 32'h13000000;
	16'h3a4 : data <= 32'hb3f12000;
	16'h3a5 : data <= 32'h13021200;
	16'h3a6 : data <= 32'h93022000;
	16'h3a7 : data <= 32'he31e52fc;
	16'h3a8 : data <= 32'hb70e0f00;
	16'h3a9 : data <= 32'h938efe00;
	16'h3aa : data <= 32'h130e1005;
	16'h3ab : data <= 32'h6384d101;
	16'h3ac : data <= 32'h6f60503a;
	16'h3ad : data <= 32'h13020000;
	16'h3ae : data <= 32'h37110f0f;
	16'h3af : data <= 32'h1301f1f0;
	16'h3b0 : data <= 32'h13000000;
	16'h3b1 : data <= 32'hb70001ff;
	16'h3b2 : data <= 32'h938000f0;
	16'h3b3 : data <= 32'hb3f12000;
	16'h3b4 : data <= 32'h13021200;
	16'h3b5 : data <= 32'h93022000;
	16'h3b6 : data <= 32'he31052fe;
	16'h3b7 : data <= 32'hb71e000f;
	16'h3b8 : data <= 32'h938e0ef0;
	16'h3b9 : data <= 32'h130e2005;
	16'h3ba : data <= 32'h6384d101;
	16'h3bb : data <= 32'h6f609036;
	16'h3bc : data <= 32'h13020000;
	16'h3bd : data <= 32'h37f1f0f0;
	16'h3be : data <= 32'h1301010f;
	16'h3bf : data <= 32'h13000000;
	16'h3c0 : data <= 32'hb710f00f;
	16'h3c1 : data <= 32'h938000ff;
	16'h3c2 : data <= 32'h13000000;
	16'h3c3 : data <= 32'hb3f12000;
	16'h3c4 : data <= 32'h13021200;
	16'h3c5 : data <= 32'h93022000;
	16'h3c6 : data <= 32'he31e52fc;
	16'h3c7 : data <= 32'hb70ef000;
	16'h3c8 : data <= 32'h938e0e0f;
	16'h3c9 : data <= 32'h130e3005;
	16'h3ca : data <= 32'h6384d101;
	16'h3cb : data <= 32'h6f609032;
	16'h3cc : data <= 32'h13020000;
	16'h3cd : data <= 32'h37110f0f;
	16'h3ce : data <= 32'h1301f1f0;
	16'h3cf : data <= 32'h13000000;
	16'h3d0 : data <= 32'h13000000;
	16'h3d1 : data <= 32'hb700ff00;
	16'h3d2 : data <= 32'h9380f00f;
	16'h3d3 : data <= 32'hb3f12000;
	16'h3d4 : data <= 32'h13021200;
	16'h3d5 : data <= 32'h93022000;
	16'h3d6 : data <= 32'he31e52fc;
	16'h3d7 : data <= 32'hb70e0f00;
	16'h3d8 : data <= 32'h938efe00;
	16'h3d9 : data <= 32'h130e4005;
	16'h3da : data <= 32'h6384d101;
	16'h3db : data <= 32'h6f60902e;
	16'h3dc : data <= 32'hb70001ff;
	16'h3dd : data <= 32'h938000f0;
	16'h3de : data <= 32'h33711000;
	16'h3df : data <= 32'h930e0000;
	16'h3e0 : data <= 32'h130e5005;
	16'h3e1 : data <= 32'h6304d101;
	16'h3e2 : data <= 32'h6f60d02c;
	16'h3e3 : data <= 32'hb700ff00;
	16'h3e4 : data <= 32'h9380f00f;
	16'h3e5 : data <= 32'h33f10000;
	16'h3e6 : data <= 32'h930e0000;
	16'h3e7 : data <= 32'h130e6005;
	16'h3e8 : data <= 32'h6304d101;
	16'h3e9 : data <= 32'h6f60102b;
	16'h3ea : data <= 32'hb3700000;
	16'h3eb : data <= 32'h930e0000;
	16'h3ec : data <= 32'h130e7005;
	16'h3ed : data <= 32'h6384d001;
	16'h3ee : data <= 32'h6f60d029;
	16'h3ef : data <= 32'hb7101111;
	16'h3f0 : data <= 32'h93801011;
	16'h3f1 : data <= 32'h37212222;
	16'h3f2 : data <= 32'h13012122;
	16'h3f3 : data <= 32'h33f02000;
	16'h3f4 : data <= 32'h930e0000;
	16'h3f5 : data <= 32'h130e8005;
	16'h3f6 : data <= 32'h6304d001;
	16'h3f7 : data <= 32'h6f609027;
	16'h3f8 : data <= 32'hb70001ff;
	16'h3f9 : data <= 32'h938000f0;
	16'h3fa : data <= 32'h93f1f0f0;
	16'h3fb : data <= 32'hb70e01ff;
	16'h3fc : data <= 32'h938e0ef0;
	16'h3fd : data <= 32'h130e9005;
	16'h3fe : data <= 32'h6384d101;
	16'h3ff : data <= 32'h6f609025;
	16'h400 : data <= 32'hb710f00f;
	16'h401 : data <= 32'h938000ff;
	16'h402 : data <= 32'h93f1000f;
	16'h403 : data <= 32'h930e000f;
	16'h404 : data <= 32'h130ea005;
	16'h405 : data <= 32'h6384d101;
	16'h406 : data <= 32'h6f60d023;
	16'h407 : data <= 32'hb700ff00;
	16'h408 : data <= 32'h9380f00f;
	16'h409 : data <= 32'h93f1f070;
	16'h40a : data <= 32'h930ef000;
	16'h40b : data <= 32'h130eb005;
	16'h40c : data <= 32'h6384d101;
	16'h40d : data <= 32'h6f601022;
	16'h40e : data <= 32'hb7f00ff0;
	16'h40f : data <= 32'h9380f000;
	16'h410 : data <= 32'h93f1000f;
	16'h411 : data <= 32'h930e0000;
	16'h412 : data <= 32'h130ec005;
	16'h413 : data <= 32'h6384d101;
	16'h414 : data <= 32'h6f605020;
	16'h415 : data <= 32'hb70001ff;
	16'h416 : data <= 32'h938000f0;
	16'h417 : data <= 32'h93f0000f;
	16'h418 : data <= 32'h930e0000;
	16'h419 : data <= 32'h130ed005;
	16'h41a : data <= 32'h6384d001;
	16'h41b : data <= 32'h6f60901e;
	16'h41c : data <= 32'h13020000;
	16'h41d : data <= 32'hb710f00f;
	16'h41e : data <= 32'h938000ff;
	16'h41f : data <= 32'h93f1f070;
	16'h420 : data <= 32'h13830100;
	16'h421 : data <= 32'h13021200;
	16'h422 : data <= 32'h93022000;
	16'h423 : data <= 32'he31452fe;
	16'h424 : data <= 32'h930e0070;
	16'h425 : data <= 32'h130ee005;
	16'h426 : data <= 32'h6304d301;
	16'h427 : data <= 32'h6f60901b;
	16'h428 : data <= 32'h13020000;
	16'h429 : data <= 32'hb700ff00;
	16'h42a : data <= 32'h9380f00f;
	16'h42b : data <= 32'h93f1000f;
	16'h42c : data <= 32'h13000000;
	16'h42d : data <= 32'h13830100;
	16'h42e : data <= 32'h13021200;
	16'h42f : data <= 32'h93022000;
	16'h430 : data <= 32'he31252fe;
	16'h431 : data <= 32'h930e000f;
	16'h432 : data <= 32'h130ef005;
	16'h433 : data <= 32'h6304d301;
	16'h434 : data <= 32'h6f605018;
	16'h435 : data <= 32'h13020000;
	16'h436 : data <= 32'hb7f00ff0;
	16'h437 : data <= 32'h9380f000;
	16'h438 : data <= 32'h93f1f0f0;
	16'h439 : data <= 32'h13000000;
	16'h43a : data <= 32'h13000000;
	16'h43b : data <= 32'h13830100;
	16'h43c : data <= 32'h13021200;
	16'h43d : data <= 32'h93022000;
	16'h43e : data <= 32'he31052fe;
	16'h43f : data <= 32'hb7fe0ff0;
	16'h440 : data <= 32'h938efe00;
	16'h441 : data <= 32'h130e0006;
	16'h442 : data <= 32'h6304d301;
	16'h443 : data <= 32'h6f609014;
	16'h444 : data <= 32'h13020000;
	16'h445 : data <= 32'hb710f00f;
	16'h446 : data <= 32'h938000ff;
	16'h447 : data <= 32'h93f1f070;
	16'h448 : data <= 32'h13021200;
	16'h449 : data <= 32'h93022000;
	16'h44a : data <= 32'he31652fe;
	16'h44b : data <= 32'h930e0070;
	16'h44c : data <= 32'h130e1006;
	16'h44d : data <= 32'h6384d101;
	16'h44e : data <= 32'h6f60d011;
	16'h44f : data <= 32'h13020000;
	16'h450 : data <= 32'hb700ff00;
	16'h451 : data <= 32'h9380f00f;
	16'h452 : data <= 32'h13000000;
	16'h453 : data <= 32'h93f1000f;
	16'h454 : data <= 32'h13021200;
	16'h455 : data <= 32'h93022000;
	16'h456 : data <= 32'he31452fe;
	16'h457 : data <= 32'h930e000f;
	16'h458 : data <= 32'h130e2006;
	16'h459 : data <= 32'h6384d101;
	16'h45a : data <= 32'h6f60d00e;
	16'h45b : data <= 32'h13020000;
	16'h45c : data <= 32'hb7f00ff0;
	16'h45d : data <= 32'h9380f000;
	16'h45e : data <= 32'h13000000;
	16'h45f : data <= 32'h13000000;
	16'h460 : data <= 32'h93f1f070;
	16'h461 : data <= 32'h13021200;
	16'h462 : data <= 32'h93022000;
	16'h463 : data <= 32'he31252fe;
	16'h464 : data <= 32'h930ef000;
	16'h465 : data <= 32'h130e3006;
	16'h466 : data <= 32'h6384d101;
	16'h467 : data <= 32'h6f60900b;
	16'h468 : data <= 32'h9370000f;
	16'h469 : data <= 32'h930e0000;
	16'h46a : data <= 32'h130e4006;
	16'h46b : data <= 32'h6384d001;
	16'h46c : data <= 32'h6f60500a;
	16'h46d : data <= 32'hb700ff00;
	16'h46e : data <= 32'h9380f00f;
	16'h46f : data <= 32'h13f0f070;
	16'h470 : data <= 32'h930e0000;
	16'h471 : data <= 32'h130e5006;
	16'h472 : data <= 32'h6304d001;
	16'h473 : data <= 32'h6f609008;
	16'h474 : data <= 32'h17250000;
	16'h475 : data <= 32'h1305c571;
	16'h476 : data <= 32'hef054000;
	16'h477 : data <= 32'h3305b540;
	16'h478 : data <= 32'hb72e0000;
	16'h479 : data <= 32'h938e0e71;
	16'h47a : data <= 32'h130e6006;
	16'h47b : data <= 32'h6304d501;
	16'h47c : data <= 32'h6f605006;
	16'h47d : data <= 32'h13000000;
	16'h47e : data <= 32'h17e5ffff;
	16'h47f : data <= 32'h1305c58f;
	16'h480 : data <= 32'hef054000;
	16'h481 : data <= 32'h3305b540;
	16'h482 : data <= 32'hb7eeffff;
	16'h483 : data <= 32'h938e0e8f;
	16'h484 : data <= 32'h130e7006;
	16'h485 : data <= 32'h6304d501;
	16'h486 : data <= 32'h6f60d003;
	16'h487 : data <= 32'h130e8006;
	16'h488 : data <= 32'h93000000;
	16'h489 : data <= 32'h13010000;
	16'h48a : data <= 32'h63882000;
	16'h48b : data <= 32'h6304c001;
	16'h48c : data <= 32'h6f605002;
	16'h48d : data <= 32'h6318c001;
	16'h48e : data <= 32'he38e20fe;
	16'h48f : data <= 32'h6304c001;
	16'h490 : data <= 32'h6f605001;
	16'h491 : data <= 32'h130e9006;
	16'h492 : data <= 32'h93001000;
	16'h493 : data <= 32'h13011000;
	16'h494 : data <= 32'h63882000;
	16'h495 : data <= 32'h6304c001;
	16'h496 : data <= 32'h6f60c07f;
	16'h497 : data <= 32'h6318c001;
	16'h498 : data <= 32'he38e20fe;
	16'h499 : data <= 32'h6304c001;
	16'h49a : data <= 32'h6f60c07e;
	16'h49b : data <= 32'h130ea006;
	16'h49c : data <= 32'h9300f0ff;
	16'h49d : data <= 32'h1301f0ff;
	16'h49e : data <= 32'h63882000;
	16'h49f : data <= 32'h6304c001;
	16'h4a0 : data <= 32'h6f60407d;
	16'h4a1 : data <= 32'h6318c001;
	16'h4a2 : data <= 32'he38e20fe;
	16'h4a3 : data <= 32'h6304c001;
	16'h4a4 : data <= 32'h6f60407c;
	16'h4a5 : data <= 32'h130eb006;
	16'h4a6 : data <= 32'h93000000;
	16'h4a7 : data <= 32'h13011000;
	16'h4a8 : data <= 32'h63842000;
	16'h4a9 : data <= 32'h6316c001;
	16'h4aa : data <= 32'h6304c001;
	16'h4ab : data <= 32'h6f60807a;
	16'h4ac : data <= 32'he38c20fe;
	16'h4ad : data <= 32'h130ec006;
	16'h4ae : data <= 32'h93001000;
	16'h4af : data <= 32'h13010000;
	16'h4b0 : data <= 32'h63842000;
	16'h4b1 : data <= 32'h6316c001;
	16'h4b2 : data <= 32'h6304c001;
	16'h4b3 : data <= 32'h6f608078;
	16'h4b4 : data <= 32'he38c20fe;
	16'h4b5 : data <= 32'h130ed006;
	16'h4b6 : data <= 32'h9300f0ff;
	16'h4b7 : data <= 32'h13011000;
	16'h4b8 : data <= 32'h63842000;
	16'h4b9 : data <= 32'h6316c001;
	16'h4ba : data <= 32'h6304c001;
	16'h4bb : data <= 32'h6f608076;
	16'h4bc : data <= 32'he38c20fe;
	16'h4bd : data <= 32'h130ee006;
	16'h4be : data <= 32'h93001000;
	16'h4bf : data <= 32'h1301f0ff;
	16'h4c0 : data <= 32'h63842000;
	16'h4c1 : data <= 32'h6316c001;
	16'h4c2 : data <= 32'h6304c001;
	16'h4c3 : data <= 32'h6f608074;
	16'h4c4 : data <= 32'he38c20fe;
	16'h4c5 : data <= 32'h130ef006;
	16'h4c6 : data <= 32'h13020000;
	16'h4c7 : data <= 32'h93000000;
	16'h4c8 : data <= 32'h1301f0ff;
	16'h4c9 : data <= 32'h63942000;
	16'h4ca : data <= 32'h6f60c072;
	16'h4cb : data <= 32'h13021200;
	16'h4cc : data <= 32'h93022000;
	16'h4cd : data <= 32'he31452fe;
	16'h4ce : data <= 32'h130e0007;
	16'h4cf : data <= 32'h13020000;
	16'h4d0 : data <= 32'h93000000;
	16'h4d1 : data <= 32'h1301f0ff;
	16'h4d2 : data <= 32'h13000000;
	16'h4d3 : data <= 32'h63942000;
	16'h4d4 : data <= 32'h6f604070;
	16'h4d5 : data <= 32'h13021200;
	16'h4d6 : data <= 32'h93022000;
	16'h4d7 : data <= 32'he31252fe;
	16'h4d8 : data <= 32'h130e1007;
	16'h4d9 : data <= 32'h13020000;
	16'h4da : data <= 32'h93000000;
	16'h4db : data <= 32'h1301f0ff;
	16'h4dc : data <= 32'h13000000;
	16'h4dd : data <= 32'h13000000;
	16'h4de : data <= 32'h63942000;
	16'h4df : data <= 32'h6f60806d;
	16'h4e0 : data <= 32'h13021200;
	16'h4e1 : data <= 32'h93022000;
	16'h4e2 : data <= 32'he31052fe;
	16'h4e3 : data <= 32'h130e2007;
	16'h4e4 : data <= 32'h13020000;
	16'h4e5 : data <= 32'h93000000;
	16'h4e6 : data <= 32'h13000000;
	16'h4e7 : data <= 32'h1301f0ff;
	16'h4e8 : data <= 32'h63942000;
	16'h4e9 : data <= 32'h6f60006b;
	16'h4ea : data <= 32'h13021200;
	16'h4eb : data <= 32'h93022000;
	16'h4ec : data <= 32'he31252fe;
	16'h4ed : data <= 32'h130e3007;
	16'h4ee : data <= 32'h13020000;
	16'h4ef : data <= 32'h93000000;
	16'h4f0 : data <= 32'h13000000;
	16'h4f1 : data <= 32'h1301f0ff;
	16'h4f2 : data <= 32'h13000000;
	16'h4f3 : data <= 32'h63942000;
	16'h4f4 : data <= 32'h6f604068;
	16'h4f5 : data <= 32'h13021200;
	16'h4f6 : data <= 32'h93022000;
	16'h4f7 : data <= 32'he31052fe;
	16'h4f8 : data <= 32'h130e4007;
	16'h4f9 : data <= 32'h13020000;
	16'h4fa : data <= 32'h93000000;
	16'h4fb : data <= 32'h13000000;
	16'h4fc : data <= 32'h13000000;
	16'h4fd : data <= 32'h1301f0ff;
	16'h4fe : data <= 32'h63942000;
	16'h4ff : data <= 32'h6f608065;
	16'h500 : data <= 32'h13021200;
	16'h501 : data <= 32'h93022000;
	16'h502 : data <= 32'he31052fe;
	16'h503 : data <= 32'h130e5007;
	16'h504 : data <= 32'h13020000;
	16'h505 : data <= 32'h93000000;
	16'h506 : data <= 32'h1301f0ff;
	16'h507 : data <= 32'h63942000;
	16'h508 : data <= 32'h6f604063;
	16'h509 : data <= 32'h13021200;
	16'h50a : data <= 32'h93022000;
	16'h50b : data <= 32'he31452fe;
	16'h50c : data <= 32'h130e6007;
	16'h50d : data <= 32'h13020000;
	16'h50e : data <= 32'h93000000;
	16'h50f : data <= 32'h1301f0ff;
	16'h510 : data <= 32'h13000000;
	16'h511 : data <= 32'h63942000;
	16'h512 : data <= 32'h6f60c060;
	16'h513 : data <= 32'h13021200;
	16'h514 : data <= 32'h93022000;
	16'h515 : data <= 32'he31252fe;
	16'h516 : data <= 32'h130e7007;
	16'h517 : data <= 32'h13020000;
	16'h518 : data <= 32'h93000000;
	16'h519 : data <= 32'h1301f0ff;
	16'h51a : data <= 32'h13000000;
	16'h51b : data <= 32'h13000000;
	16'h51c : data <= 32'h63942000;
	16'h51d : data <= 32'h6f60005e;
	16'h51e : data <= 32'h13021200;
	16'h51f : data <= 32'h93022000;
	16'h520 : data <= 32'he31052fe;
	16'h521 : data <= 32'h130e8007;
	16'h522 : data <= 32'h13020000;
	16'h523 : data <= 32'h93000000;
	16'h524 : data <= 32'h13000000;
	16'h525 : data <= 32'h1301f0ff;
	16'h526 : data <= 32'h63942000;
	16'h527 : data <= 32'h6f60805b;
	16'h528 : data <= 32'h13021200;
	16'h529 : data <= 32'h93022000;
	16'h52a : data <= 32'he31252fe;
	16'h52b : data <= 32'h130e9007;
	16'h52c : data <= 32'h13020000;
	16'h52d : data <= 32'h93000000;
	16'h52e : data <= 32'h13000000;
	16'h52f : data <= 32'h1301f0ff;
	16'h530 : data <= 32'h13000000;
	16'h531 : data <= 32'h63942000;
	16'h532 : data <= 32'h6f60c058;
	16'h533 : data <= 32'h13021200;
	16'h534 : data <= 32'h93022000;
	16'h535 : data <= 32'he31052fe;
	16'h536 : data <= 32'h130ea007;
	16'h537 : data <= 32'h13020000;
	16'h538 : data <= 32'h93000000;
	16'h539 : data <= 32'h13000000;
	16'h53a : data <= 32'h13000000;
	16'h53b : data <= 32'h1301f0ff;
	16'h53c : data <= 32'h63942000;
	16'h53d : data <= 32'h6f600056;
	16'h53e : data <= 32'h13021200;
	16'h53f : data <= 32'h93022000;
	16'h540 : data <= 32'he31052fe;
	16'h541 : data <= 32'h93001000;
	16'h542 : data <= 32'h630a0000;
	16'h543 : data <= 32'h93801000;
	16'h544 : data <= 32'h93801000;
	16'h545 : data <= 32'h93801000;
	16'h546 : data <= 32'h93801000;
	16'h547 : data <= 32'h93801000;
	16'h548 : data <= 32'h93801000;
	16'h549 : data <= 32'h930e3000;
	16'h54a : data <= 32'h130eb007;
	16'h54b : data <= 32'h6384d001;
	16'h54c : data <= 32'h6f604052;
	16'h54d : data <= 32'h130ec007;
	16'h54e : data <= 32'h93000000;
	16'h54f : data <= 32'h13010000;
	16'h550 : data <= 32'h63d82000;
	16'h551 : data <= 32'h6304c001;
	16'h552 : data <= 32'h6f60c050;
	16'h553 : data <= 32'h6318c001;
	16'h554 : data <= 32'he3de20fe;
	16'h555 : data <= 32'h6304c001;
	16'h556 : data <= 32'h6f60c04f;
	16'h557 : data <= 32'h130ed007;
	16'h558 : data <= 32'h93001000;
	16'h559 : data <= 32'h13011000;
	16'h55a : data <= 32'h63d82000;
	16'h55b : data <= 32'h6304c001;
	16'h55c : data <= 32'h6f60404e;
	16'h55d : data <= 32'h6318c001;
	16'h55e : data <= 32'he3de20fe;
	16'h55f : data <= 32'h6304c001;
	16'h560 : data <= 32'h6f60404d;
	16'h561 : data <= 32'h130ee007;
	16'h562 : data <= 32'h9300f0ff;
	16'h563 : data <= 32'h1301f0ff;
	16'h564 : data <= 32'h63d82000;
	16'h565 : data <= 32'h6304c001;
	16'h566 : data <= 32'h6f60c04b;
	16'h567 : data <= 32'h6318c001;
	16'h568 : data <= 32'he3de20fe;
	16'h569 : data <= 32'h6304c001;
	16'h56a : data <= 32'h6f60c04a;
	16'h56b : data <= 32'h130ef007;
	16'h56c : data <= 32'h93001000;
	16'h56d : data <= 32'h13010000;
	16'h56e : data <= 32'h63d82000;
	16'h56f : data <= 32'h6304c001;
	16'h570 : data <= 32'h6f604049;
	16'h571 : data <= 32'h6318c001;
	16'h572 : data <= 32'he3de20fe;
	16'h573 : data <= 32'h6304c001;
	16'h574 : data <= 32'h6f604048;
	16'h575 : data <= 32'h130e0008;
	16'h576 : data <= 32'h93001000;
	16'h577 : data <= 32'h1301f0ff;
	16'h578 : data <= 32'h63d82000;
	16'h579 : data <= 32'h6304c001;
	16'h57a : data <= 32'h6f60c046;
	16'h57b : data <= 32'h6318c001;
	16'h57c : data <= 32'he3de20fe;
	16'h57d : data <= 32'h6304c001;
	16'h57e : data <= 32'h6f60c045;
	16'h57f : data <= 32'h130e1008;
	16'h580 : data <= 32'h9300f0ff;
	16'h581 : data <= 32'h1301e0ff;
	16'h582 : data <= 32'h63d82000;
	16'h583 : data <= 32'h6304c001;
	16'h584 : data <= 32'h6f604044;
	16'h585 : data <= 32'h6318c001;
	16'h586 : data <= 32'he3de20fe;
	16'h587 : data <= 32'h6304c001;
	16'h588 : data <= 32'h6f604043;
	16'h589 : data <= 32'h130e2008;
	16'h58a : data <= 32'h93000000;
	16'h58b : data <= 32'h13011000;
	16'h58c : data <= 32'h63d42000;
	16'h58d : data <= 32'h6316c001;
	16'h58e : data <= 32'h6304c001;
	16'h58f : data <= 32'h6f608041;
	16'h590 : data <= 32'he3dc20fe;
	16'h591 : data <= 32'h130e3008;
	16'h592 : data <= 32'h9300f0ff;
	16'h593 : data <= 32'h13011000;
	16'h594 : data <= 32'h63d42000;
	16'h595 : data <= 32'h6316c001;
	16'h596 : data <= 32'h6304c001;
	16'h597 : data <= 32'h6f60803f;
	16'h598 : data <= 32'he3dc20fe;
	16'h599 : data <= 32'h130e4008;
	16'h59a : data <= 32'h9300e0ff;
	16'h59b : data <= 32'h1301f0ff;
	16'h59c : data <= 32'h63d42000;
	16'h59d : data <= 32'h6316c001;
	16'h59e : data <= 32'h6304c001;
	16'h59f : data <= 32'h6f60803d;
	16'h5a0 : data <= 32'he3dc20fe;
	16'h5a1 : data <= 32'h130e5008;
	16'h5a2 : data <= 32'h9300e0ff;
	16'h5a3 : data <= 32'h13011000;
	16'h5a4 : data <= 32'h63d42000;
	16'h5a5 : data <= 32'h6316c001;
	16'h5a6 : data <= 32'h6304c001;
	16'h5a7 : data <= 32'h6f60803b;
	16'h5a8 : data <= 32'he3dc20fe;
	16'h5a9 : data <= 32'h130e6008;
	16'h5aa : data <= 32'h13020000;
	16'h5ab : data <= 32'h9300f0ff;
	16'h5ac : data <= 32'h13010000;
	16'h5ad : data <= 32'h63c42000;
	16'h5ae : data <= 32'h6f60c039;
	16'h5af : data <= 32'h13021200;
	16'h5b0 : data <= 32'h93022000;
	16'h5b1 : data <= 32'he31452fe;
	16'h5b2 : data <= 32'h130e7008;
	16'h5b3 : data <= 32'h13020000;
	16'h5b4 : data <= 32'h9300f0ff;
	16'h5b5 : data <= 32'h13010000;
	16'h5b6 : data <= 32'h13000000;
	16'h5b7 : data <= 32'h63c42000;
	16'h5b8 : data <= 32'h6f604037;
	16'h5b9 : data <= 32'h13021200;
	16'h5ba : data <= 32'h93022000;
	16'h5bb : data <= 32'he31252fe;
	16'h5bc : data <= 32'h130e8008;
	16'h5bd : data <= 32'h13020000;
	16'h5be : data <= 32'h9300f0ff;
	16'h5bf : data <= 32'h13010000;
	16'h5c0 : data <= 32'h13000000;
	16'h5c1 : data <= 32'h13000000;
	16'h5c2 : data <= 32'h63c42000;
	16'h5c3 : data <= 32'h6f608034;
	16'h5c4 : data <= 32'h13021200;
	16'h5c5 : data <= 32'h93022000;
	16'h5c6 : data <= 32'he31052fe;
	16'h5c7 : data <= 32'h130e9008;
	16'h5c8 : data <= 32'h13020000;
	16'h5c9 : data <= 32'h9300f0ff;
	16'h5ca : data <= 32'h13000000;
	16'h5cb : data <= 32'h13010000;
	16'h5cc : data <= 32'h63c42000;
	16'h5cd : data <= 32'h6f600032;
	16'h5ce : data <= 32'h13021200;
	16'h5cf : data <= 32'h93022000;
	16'h5d0 : data <= 32'he31252fe;
	16'h5d1 : data <= 32'h130ea008;
	16'h5d2 : data <= 32'h13020000;
	16'h5d3 : data <= 32'h9300f0ff;
	16'h5d4 : data <= 32'h13000000;
	16'h5d5 : data <= 32'h13010000;
	16'h5d6 : data <= 32'h13000000;
	16'h5d7 : data <= 32'h63c42000;
	16'h5d8 : data <= 32'h6f60402f;
	16'h5d9 : data <= 32'h13021200;
	16'h5da : data <= 32'h93022000;
	16'h5db : data <= 32'he31052fe;
	16'h5dc : data <= 32'h130eb008;
	16'h5dd : data <= 32'h13020000;
	16'h5de : data <= 32'h9300f0ff;
	16'h5df : data <= 32'h13000000;
	16'h5e0 : data <= 32'h13000000;
	16'h5e1 : data <= 32'h13010000;
	16'h5e2 : data <= 32'h63c42000;
	16'h5e3 : data <= 32'h6f60802c;
	16'h5e4 : data <= 32'h13021200;
	16'h5e5 : data <= 32'h93022000;
	16'h5e6 : data <= 32'he31052fe;
	16'h5e7 : data <= 32'h130ec008;
	16'h5e8 : data <= 32'h13020000;
	16'h5e9 : data <= 32'h9300f0ff;
	16'h5ea : data <= 32'h13010000;
	16'h5eb : data <= 32'h63c42000;
	16'h5ec : data <= 32'h6f60402a;
	16'h5ed : data <= 32'h13021200;
	16'h5ee : data <= 32'h93022000;
	16'h5ef : data <= 32'he31452fe;
	16'h5f0 : data <= 32'h130ed008;
	16'h5f1 : data <= 32'h13020000;
	16'h5f2 : data <= 32'h9300f0ff;
	16'h5f3 : data <= 32'h13010000;
	16'h5f4 : data <= 32'h13000000;
	16'h5f5 : data <= 32'h63c42000;
	16'h5f6 : data <= 32'h6f60c027;
	16'h5f7 : data <= 32'h13021200;
	16'h5f8 : data <= 32'h93022000;
	16'h5f9 : data <= 32'he31252fe;
	16'h5fa : data <= 32'h130ee008;
	16'h5fb : data <= 32'h13020000;
	16'h5fc : data <= 32'h9300f0ff;
	16'h5fd : data <= 32'h13010000;
	16'h5fe : data <= 32'h13000000;
	16'h5ff : data <= 32'h13000000;
	16'h600 : data <= 32'h63c42000;
	16'h601 : data <= 32'h6f600025;
	16'h602 : data <= 32'h13021200;
	16'h603 : data <= 32'h93022000;
	16'h604 : data <= 32'he31052fe;
	16'h605 : data <= 32'h130ef008;
	16'h606 : data <= 32'h13020000;
	16'h607 : data <= 32'h9300f0ff;
	16'h608 : data <= 32'h13000000;
	16'h609 : data <= 32'h13010000;
	16'h60a : data <= 32'h63c42000;
	16'h60b : data <= 32'h6f608022;
	16'h60c : data <= 32'h13021200;
	16'h60d : data <= 32'h93022000;
	16'h60e : data <= 32'he31252fe;
	16'h60f : data <= 32'h130e0009;
	16'h610 : data <= 32'h13020000;
	16'h611 : data <= 32'h9300f0ff;
	16'h612 : data <= 32'h13000000;
	16'h613 : data <= 32'h13010000;
	16'h614 : data <= 32'h13000000;
	16'h615 : data <= 32'h63c42000;
	16'h616 : data <= 32'h6f60c01f;
	16'h617 : data <= 32'h13021200;
	16'h618 : data <= 32'h93022000;
	16'h619 : data <= 32'he31052fe;
	16'h61a : data <= 32'h130e1009;
	16'h61b : data <= 32'h13020000;
	16'h61c : data <= 32'h9300f0ff;
	16'h61d : data <= 32'h13000000;
	16'h61e : data <= 32'h13000000;
	16'h61f : data <= 32'h13010000;
	16'h620 : data <= 32'h63c42000;
	16'h621 : data <= 32'h6f60001d;
	16'h622 : data <= 32'h13021200;
	16'h623 : data <= 32'h93022000;
	16'h624 : data <= 32'he31052fe;
	16'h625 : data <= 32'h93001000;
	16'h626 : data <= 32'h63da0000;
	16'h627 : data <= 32'h93801000;
	16'h628 : data <= 32'h93801000;
	16'h629 : data <= 32'h93801000;
	16'h62a : data <= 32'h93801000;
	16'h62b : data <= 32'h93801000;
	16'h62c : data <= 32'h93801000;
	16'h62d : data <= 32'h930e3000;
	16'h62e : data <= 32'h130e2009;
	16'h62f : data <= 32'h6384d001;
	16'h630 : data <= 32'h6f604019;
	16'h631 : data <= 32'h130e3009;
	16'h632 : data <= 32'h93000000;
	16'h633 : data <= 32'h13010000;
	16'h634 : data <= 32'h63f82000;
	16'h635 : data <= 32'h6304c001;
	16'h636 : data <= 32'h6f60c017;
	16'h637 : data <= 32'h6318c001;
	16'h638 : data <= 32'he3fe20fe;
	16'h639 : data <= 32'h6304c001;
	16'h63a : data <= 32'h6f60c016;
	16'h63b : data <= 32'h130e4009;
	16'h63c : data <= 32'h93001000;
	16'h63d : data <= 32'h13011000;
	16'h63e : data <= 32'h63f82000;
	16'h63f : data <= 32'h6304c001;
	16'h640 : data <= 32'h6f604015;
	16'h641 : data <= 32'h6318c001;
	16'h642 : data <= 32'he3fe20fe;
	16'h643 : data <= 32'h6304c001;
	16'h644 : data <= 32'h6f604014;
	16'h645 : data <= 32'h130e5009;
	16'h646 : data <= 32'h9300f0ff;
	16'h647 : data <= 32'h1301f0ff;
	16'h648 : data <= 32'h63f82000;
	16'h649 : data <= 32'h6304c001;
	16'h64a : data <= 32'h6f60c012;
	16'h64b : data <= 32'h6318c001;
	16'h64c : data <= 32'he3fe20fe;
	16'h64d : data <= 32'h6304c001;
	16'h64e : data <= 32'h6f60c011;
	16'h64f : data <= 32'h130e6009;
	16'h650 : data <= 32'h93001000;
	16'h651 : data <= 32'h13010000;
	16'h652 : data <= 32'h63f82000;
	16'h653 : data <= 32'h6304c001;
	16'h654 : data <= 32'h6f604010;
	16'h655 : data <= 32'h6318c001;
	16'h656 : data <= 32'he3fe20fe;
	16'h657 : data <= 32'h6304c001;
	16'h658 : data <= 32'h6f60400f;
	16'h659 : data <= 32'h130e7009;
	16'h65a : data <= 32'h9300f0ff;
	16'h65b : data <= 32'h1301e0ff;
	16'h65c : data <= 32'h63f82000;
	16'h65d : data <= 32'h6304c001;
	16'h65e : data <= 32'h6f60c00d;
	16'h65f : data <= 32'h6318c001;
	16'h660 : data <= 32'he3fe20fe;
	16'h661 : data <= 32'h6304c001;
	16'h662 : data <= 32'h6f60c00c;
	16'h663 : data <= 32'h130e8009;
	16'h664 : data <= 32'h9300f0ff;
	16'h665 : data <= 32'h13010000;
	16'h666 : data <= 32'h63f82000;
	16'h667 : data <= 32'h6304c001;
	16'h668 : data <= 32'h6f60400b;
	16'h669 : data <= 32'h6318c001;
	16'h66a : data <= 32'he3fe20fe;
	16'h66b : data <= 32'h6304c001;
	16'h66c : data <= 32'h6f60400a;
	16'h66d : data <= 32'h130e9009;
	16'h66e : data <= 32'h93000000;
	16'h66f : data <= 32'h13011000;
	16'h670 : data <= 32'h63f42000;
	16'h671 : data <= 32'h6316c001;
	16'h672 : data <= 32'h6304c001;
	16'h673 : data <= 32'h6f608008;
	16'h674 : data <= 32'he3fc20fe;
	16'h675 : data <= 32'h130ea009;
	16'h676 : data <= 32'h9300e0ff;
	16'h677 : data <= 32'h1301f0ff;
	16'h678 : data <= 32'h63f42000;
	16'h679 : data <= 32'h6316c001;
	16'h67a : data <= 32'h6304c001;
	16'h67b : data <= 32'h6f608006;
	16'h67c : data <= 32'he3fc20fe;
	16'h67d : data <= 32'h130eb009;
	16'h67e : data <= 32'h93000000;
	16'h67f : data <= 32'h1301f0ff;
	16'h680 : data <= 32'h63f42000;
	16'h681 : data <= 32'h6316c001;
	16'h682 : data <= 32'h6304c001;
	16'h683 : data <= 32'h6f608004;
	16'h684 : data <= 32'he3fc20fe;
	16'h685 : data <= 32'h130ec009;
	16'h686 : data <= 32'hb7000080;
	16'h687 : data <= 32'h9380f0ff;
	16'h688 : data <= 32'h37010080;
	16'h689 : data <= 32'h63f42000;
	16'h68a : data <= 32'h6316c001;
	16'h68b : data <= 32'h6304c001;
	16'h68c : data <= 32'h6f604002;
	16'h68d : data <= 32'he3fc20fe;
	16'h68e : data <= 32'h130ed009;
	16'h68f : data <= 32'h13020000;
	16'h690 : data <= 32'hb70000f0;
	16'h691 : data <= 32'h9380f0ff;
	16'h692 : data <= 32'h370100f0;
	16'h693 : data <= 32'h63e42000;
	16'h694 : data <= 32'h6f604000;
	16'h695 : data <= 32'h13021200;
	16'h696 : data <= 32'h93022000;
	16'h697 : data <= 32'he31252fe;
	16'h698 : data <= 32'h130ee009;
	16'h699 : data <= 32'h13020000;
	16'h69a : data <= 32'hb70000f0;
	16'h69b : data <= 32'h9380f0ff;
	16'h69c : data <= 32'h370100f0;
	16'h69d : data <= 32'h13000000;
	16'h69e : data <= 32'h63e42000;
	16'h69f : data <= 32'h6f50907d;
	16'h6a0 : data <= 32'h13021200;
	16'h6a1 : data <= 32'h93022000;
	16'h6a2 : data <= 32'he31052fe;
	16'h6a3 : data <= 32'h130ef009;
	16'h6a4 : data <= 32'h13020000;
	16'h6a5 : data <= 32'hb70000f0;
	16'h6a6 : data <= 32'h9380f0ff;
	16'h6a7 : data <= 32'h370100f0;
	16'h6a8 : data <= 32'h13000000;
	16'h6a9 : data <= 32'h13000000;
	16'h6aa : data <= 32'h63e42000;
	16'h6ab : data <= 32'h6f50907a;
	16'h6ac : data <= 32'h13021200;
	16'h6ad : data <= 32'h93022000;
	16'h6ae : data <= 32'he31e52fc;
	16'h6af : data <= 32'h130e000a;
	16'h6b0 : data <= 32'h13020000;
	16'h6b1 : data <= 32'hb70000f0;
	16'h6b2 : data <= 32'h9380f0ff;
	16'h6b3 : data <= 32'h13000000;
	16'h6b4 : data <= 32'h370100f0;
	16'h6b5 : data <= 32'h63e42000;
	16'h6b6 : data <= 32'h6f50d077;
	16'h6b7 : data <= 32'h13021200;
	16'h6b8 : data <= 32'h93022000;
	16'h6b9 : data <= 32'he31052fe;
	16'h6ba : data <= 32'h130e100a;
	16'h6bb : data <= 32'h13020000;
	16'h6bc : data <= 32'hb70000f0;
	16'h6bd : data <= 32'h9380f0ff;
	16'h6be : data <= 32'h13000000;
	16'h6bf : data <= 32'h370100f0;
	16'h6c0 : data <= 32'h13000000;
	16'h6c1 : data <= 32'h63e42000;
	16'h6c2 : data <= 32'h6f50d074;
	16'h6c3 : data <= 32'h13021200;
	16'h6c4 : data <= 32'h93022000;
	16'h6c5 : data <= 32'he31e52fc;
	16'h6c6 : data <= 32'h130e200a;
	16'h6c7 : data <= 32'h13020000;
	16'h6c8 : data <= 32'hb70000f0;
	16'h6c9 : data <= 32'h9380f0ff;
	16'h6ca : data <= 32'h13000000;
	16'h6cb : data <= 32'h13000000;
	16'h6cc : data <= 32'h370100f0;
	16'h6cd : data <= 32'h63e42000;
	16'h6ce : data <= 32'h6f50d071;
	16'h6cf : data <= 32'h13021200;
	16'h6d0 : data <= 32'h93022000;
	16'h6d1 : data <= 32'he31e52fc;
	16'h6d2 : data <= 32'h130e300a;
	16'h6d3 : data <= 32'h13020000;
	16'h6d4 : data <= 32'hb70000f0;
	16'h6d5 : data <= 32'h9380f0ff;
	16'h6d6 : data <= 32'h370100f0;
	16'h6d7 : data <= 32'h63e42000;
	16'h6d8 : data <= 32'h6f50506f;
	16'h6d9 : data <= 32'h13021200;
	16'h6da : data <= 32'h93022000;
	16'h6db : data <= 32'he31252fe;
	16'h6dc : data <= 32'h130e400a;
	16'h6dd : data <= 32'h13020000;
	16'h6de : data <= 32'hb70000f0;
	16'h6df : data <= 32'h9380f0ff;
	16'h6e0 : data <= 32'h370100f0;
	16'h6e1 : data <= 32'h13000000;
	16'h6e2 : data <= 32'h63e42000;
	16'h6e3 : data <= 32'h6f50906c;
	16'h6e4 : data <= 32'h13021200;
	16'h6e5 : data <= 32'h93022000;
	16'h6e6 : data <= 32'he31052fe;
	16'h6e7 : data <= 32'h130e500a;
	16'h6e8 : data <= 32'h13020000;
	16'h6e9 : data <= 32'hb70000f0;
	16'h6ea : data <= 32'h9380f0ff;
	16'h6eb : data <= 32'h370100f0;
	16'h6ec : data <= 32'h13000000;
	16'h6ed : data <= 32'h13000000;
	16'h6ee : data <= 32'h63e42000;
	16'h6ef : data <= 32'h6f509069;
	16'h6f0 : data <= 32'h13021200;
	16'h6f1 : data <= 32'h93022000;
	16'h6f2 : data <= 32'he31e52fc;
	16'h6f3 : data <= 32'h130e600a;
	16'h6f4 : data <= 32'h13020000;
	16'h6f5 : data <= 32'hb70000f0;
	16'h6f6 : data <= 32'h9380f0ff;
	16'h6f7 : data <= 32'h13000000;
	16'h6f8 : data <= 32'h370100f0;
	16'h6f9 : data <= 32'h63e42000;
	16'h6fa : data <= 32'h6f50d066;
	16'h6fb : data <= 32'h13021200;
	16'h6fc : data <= 32'h93022000;
	16'h6fd : data <= 32'he31052fe;
	16'h6fe : data <= 32'h130e700a;
	16'h6ff : data <= 32'h13020000;
	16'h700 : data <= 32'hb70000f0;
	16'h701 : data <= 32'h9380f0ff;
	16'h702 : data <= 32'h13000000;
	16'h703 : data <= 32'h370100f0;
	16'h704 : data <= 32'h13000000;
	16'h705 : data <= 32'h63e42000;
	16'h706 : data <= 32'h6f50d063;
	16'h707 : data <= 32'h13021200;
	16'h708 : data <= 32'h93022000;
	16'h709 : data <= 32'he31e52fc;
	16'h70a : data <= 32'h130e800a;
	16'h70b : data <= 32'h13020000;
	16'h70c : data <= 32'hb70000f0;
	16'h70d : data <= 32'h9380f0ff;
	16'h70e : data <= 32'h13000000;
	16'h70f : data <= 32'h13000000;
	16'h710 : data <= 32'h370100f0;
	16'h711 : data <= 32'h63e42000;
	16'h712 : data <= 32'h6f50d060;
	16'h713 : data <= 32'h13021200;
	16'h714 : data <= 32'h93022000;
	16'h715 : data <= 32'he31e52fc;
	16'h716 : data <= 32'h93001000;
	16'h717 : data <= 32'h63fa0000;
	16'h718 : data <= 32'h93801000;
	16'h719 : data <= 32'h93801000;
	16'h71a : data <= 32'h93801000;
	16'h71b : data <= 32'h93801000;
	16'h71c : data <= 32'h93801000;
	16'h71d : data <= 32'h93801000;
	16'h71e : data <= 32'h930e3000;
	16'h71f : data <= 32'h130e900a;
	16'h720 : data <= 32'h6384d001;
	16'h721 : data <= 32'h6f50105d;
	16'h722 : data <= 32'h130ea00a;
	16'h723 : data <= 32'h93000000;
	16'h724 : data <= 32'h13011000;
	16'h725 : data <= 32'h63c82000;
	16'h726 : data <= 32'h6304c001;
	16'h727 : data <= 32'h6f50905b;
	16'h728 : data <= 32'h6318c001;
	16'h729 : data <= 32'he3ce20fe;
	16'h72a : data <= 32'h6304c001;
	16'h72b : data <= 32'h6f50905a;
	16'h72c : data <= 32'h130eb00a;
	16'h72d : data <= 32'h9300f0ff;
	16'h72e : data <= 32'h13011000;
	16'h72f : data <= 32'h63c82000;
	16'h730 : data <= 32'h6304c001;
	16'h731 : data <= 32'h6f501059;
	16'h732 : data <= 32'h6318c001;
	16'h733 : data <= 32'he3ce20fe;
	16'h734 : data <= 32'h6304c001;
	16'h735 : data <= 32'h6f501058;
	16'h736 : data <= 32'h130ec00a;
	16'h737 : data <= 32'h9300e0ff;
	16'h738 : data <= 32'h1301f0ff;
	16'h739 : data <= 32'h63c82000;
	16'h73a : data <= 32'h6304c001;
	16'h73b : data <= 32'h6f509056;
	16'h73c : data <= 32'h6318c001;
	16'h73d : data <= 32'he3ce20fe;
	16'h73e : data <= 32'h6304c001;
	16'h73f : data <= 32'h6f509055;
	16'h740 : data <= 32'h130ed00a;
	16'h741 : data <= 32'h93001000;
	16'h742 : data <= 32'h13010000;
	16'h743 : data <= 32'h63c42000;
	16'h744 : data <= 32'h6316c001;
	16'h745 : data <= 32'h6304c001;
	16'h746 : data <= 32'h6f50d053;
	16'h747 : data <= 32'he3cc20fe;
	16'h748 : data <= 32'h130ee00a;
	16'h749 : data <= 32'h93001000;
	16'h74a : data <= 32'h1301f0ff;
	16'h74b : data <= 32'h63c42000;
	16'h74c : data <= 32'h6316c001;
	16'h74d : data <= 32'h6304c001;
	16'h74e : data <= 32'h6f50d051;
	16'h74f : data <= 32'he3cc20fe;
	16'h750 : data <= 32'h130ef00a;
	16'h751 : data <= 32'h9300f0ff;
	16'h752 : data <= 32'h1301e0ff;
	16'h753 : data <= 32'h63c42000;
	16'h754 : data <= 32'h6316c001;
	16'h755 : data <= 32'h6304c001;
	16'h756 : data <= 32'h6f50d04f;
	16'h757 : data <= 32'he3cc20fe;
	16'h758 : data <= 32'h130e000b;
	16'h759 : data <= 32'h93001000;
	16'h75a : data <= 32'h1301e0ff;
	16'h75b : data <= 32'h63c42000;
	16'h75c : data <= 32'h6316c001;
	16'h75d : data <= 32'h6304c001;
	16'h75e : data <= 32'h6f50d04d;
	16'h75f : data <= 32'he3cc20fe;
	16'h760 : data <= 32'h130e100b;
	16'h761 : data <= 32'h13020000;
	16'h762 : data <= 32'h93000000;
	16'h763 : data <= 32'h1301f0ff;
	16'h764 : data <= 32'h63d42000;
	16'h765 : data <= 32'h6f50104c;
	16'h766 : data <= 32'h13021200;
	16'h767 : data <= 32'h93022000;
	16'h768 : data <= 32'he31452fe;
	16'h769 : data <= 32'h130e200b;
	16'h76a : data <= 32'h13020000;
	16'h76b : data <= 32'h93000000;
	16'h76c : data <= 32'h1301f0ff;
	16'h76d : data <= 32'h13000000;
	16'h76e : data <= 32'h63d42000;
	16'h76f : data <= 32'h6f509049;
	16'h770 : data <= 32'h13021200;
	16'h771 : data <= 32'h93022000;
	16'h772 : data <= 32'he31252fe;
	16'h773 : data <= 32'h130e300b;
	16'h774 : data <= 32'h13020000;
	16'h775 : data <= 32'h93000000;
	16'h776 : data <= 32'h1301f0ff;
	16'h777 : data <= 32'h13000000;
	16'h778 : data <= 32'h13000000;
	16'h779 : data <= 32'h63d42000;
	16'h77a : data <= 32'h6f50d046;
	16'h77b : data <= 32'h13021200;
	16'h77c : data <= 32'h93022000;
	16'h77d : data <= 32'he31052fe;
	16'h77e : data <= 32'h130e400b;
	16'h77f : data <= 32'h13020000;
	16'h780 : data <= 32'h93000000;
	16'h781 : data <= 32'h13000000;
	16'h782 : data <= 32'h1301f0ff;
	16'h783 : data <= 32'h63d42000;
	16'h784 : data <= 32'h6f505044;
	16'h785 : data <= 32'h13021200;
	16'h786 : data <= 32'h93022000;
	16'h787 : data <= 32'he31252fe;
	16'h788 : data <= 32'h130e500b;
	16'h789 : data <= 32'h13020000;
	16'h78a : data <= 32'h93000000;
	16'h78b : data <= 32'h13000000;
	16'h78c : data <= 32'h1301f0ff;
	16'h78d : data <= 32'h13000000;
	16'h78e : data <= 32'h63d42000;
	16'h78f : data <= 32'h6f509041;
	16'h790 : data <= 32'h13021200;
	16'h791 : data <= 32'h93022000;
	16'h792 : data <= 32'he31052fe;
	16'h793 : data <= 32'h130e600b;
	16'h794 : data <= 32'h13020000;
	16'h795 : data <= 32'h93000000;
	16'h796 : data <= 32'h13000000;
	16'h797 : data <= 32'h13000000;
	16'h798 : data <= 32'h1301f0ff;
	16'h799 : data <= 32'h63d42000;
	16'h79a : data <= 32'h6f50d03e;
	16'h79b : data <= 32'h13021200;
	16'h79c : data <= 32'h93022000;
	16'h79d : data <= 32'he31052fe;
	16'h79e : data <= 32'h130e700b;
	16'h79f : data <= 32'h13020000;
	16'h7a0 : data <= 32'h93000000;
	16'h7a1 : data <= 32'h1301f0ff;
	16'h7a2 : data <= 32'h63d42000;
	16'h7a3 : data <= 32'h6f50903c;
	16'h7a4 : data <= 32'h13021200;
	16'h7a5 : data <= 32'h93022000;
	16'h7a6 : data <= 32'he31452fe;
	16'h7a7 : data <= 32'h130e800b;
	16'h7a8 : data <= 32'h13020000;
	16'h7a9 : data <= 32'h93000000;
	16'h7aa : data <= 32'h1301f0ff;
	16'h7ab : data <= 32'h13000000;
	16'h7ac : data <= 32'h63d42000;
	16'h7ad : data <= 32'h6f50103a;
	16'h7ae : data <= 32'h13021200;
	16'h7af : data <= 32'h93022000;
	16'h7b0 : data <= 32'he31252fe;
	16'h7b1 : data <= 32'h130e900b;
	16'h7b2 : data <= 32'h13020000;
	16'h7b3 : data <= 32'h93000000;
	16'h7b4 : data <= 32'h1301f0ff;
	16'h7b5 : data <= 32'h13000000;
	16'h7b6 : data <= 32'h13000000;
	16'h7b7 : data <= 32'h63d42000;
	16'h7b8 : data <= 32'h6f505037;
	16'h7b9 : data <= 32'h13021200;
	16'h7ba : data <= 32'h93022000;
	16'h7bb : data <= 32'he31052fe;
	16'h7bc : data <= 32'h130ea00b;
	16'h7bd : data <= 32'h13020000;
	16'h7be : data <= 32'h93000000;
	16'h7bf : data <= 32'h13000000;
	16'h7c0 : data <= 32'h1301f0ff;
	16'h7c1 : data <= 32'h63d42000;
	16'h7c2 : data <= 32'h6f50d034;
	16'h7c3 : data <= 32'h13021200;
	16'h7c4 : data <= 32'h93022000;
	16'h7c5 : data <= 32'he31252fe;
	16'h7c6 : data <= 32'h130eb00b;
	16'h7c7 : data <= 32'h13020000;
	16'h7c8 : data <= 32'h93000000;
	16'h7c9 : data <= 32'h13000000;
	16'h7ca : data <= 32'h1301f0ff;
	16'h7cb : data <= 32'h13000000;
	16'h7cc : data <= 32'h63d42000;
	16'h7cd : data <= 32'h6f501032;
	16'h7ce : data <= 32'h13021200;
	16'h7cf : data <= 32'h93022000;
	16'h7d0 : data <= 32'he31052fe;
	16'h7d1 : data <= 32'h130ec00b;
	16'h7d2 : data <= 32'h13020000;
	16'h7d3 : data <= 32'h93000000;
	16'h7d4 : data <= 32'h13000000;
	16'h7d5 : data <= 32'h13000000;
	16'h7d6 : data <= 32'h1301f0ff;
	16'h7d7 : data <= 32'h63d42000;
	16'h7d8 : data <= 32'h6f50502f;
	16'h7d9 : data <= 32'h13021200;
	16'h7da : data <= 32'h93022000;
	16'h7db : data <= 32'he31052fe;
	16'h7dc : data <= 32'h93001000;
	16'h7dd : data <= 32'h634a1000;
	16'h7de : data <= 32'h93801000;
	16'h7df : data <= 32'h93801000;
	16'h7e0 : data <= 32'h93801000;
	16'h7e1 : data <= 32'h93801000;
	16'h7e2 : data <= 32'h93801000;
	16'h7e3 : data <= 32'h93801000;
	16'h7e4 : data <= 32'h930e3000;
	16'h7e5 : data <= 32'h130ed00b;
	16'h7e6 : data <= 32'h6384d001;
	16'h7e7 : data <= 32'h6f50902b;
	16'h7e8 : data <= 32'h130ee00b;
	16'h7e9 : data <= 32'h93000000;
	16'h7ea : data <= 32'h13011000;
	16'h7eb : data <= 32'h63e82000;
	16'h7ec : data <= 32'h6304c001;
	16'h7ed : data <= 32'h6f50102a;
	16'h7ee : data <= 32'h6318c001;
	16'h7ef : data <= 32'he3ee20fe;
	16'h7f0 : data <= 32'h6304c001;
	16'h7f1 : data <= 32'h6f501029;
	16'h7f2 : data <= 32'h130ef00b;
	16'h7f3 : data <= 32'h9300e0ff;
	16'h7f4 : data <= 32'h1301f0ff;
	16'h7f5 : data <= 32'h63e82000;
	16'h7f6 : data <= 32'h6304c001;
	16'h7f7 : data <= 32'h6f509027;
	16'h7f8 : data <= 32'h6318c001;
	16'h7f9 : data <= 32'he3ee20fe;
	16'h7fa : data <= 32'h6304c001;
	16'h7fb : data <= 32'h6f509026;
	16'h7fc : data <= 32'h130e000c;
	16'h7fd : data <= 32'h93000000;
	16'h7fe : data <= 32'h1301f0ff;
	16'h7ff : data <= 32'h63e82000;
	16'h800 : data <= 32'h6304c001;
	16'h801 : data <= 32'h6f501025;
	16'h802 : data <= 32'h6318c001;
	16'h803 : data <= 32'he3ee20fe;
	16'h804 : data <= 32'h6304c001;
	16'h805 : data <= 32'h6f501024;
	16'h806 : data <= 32'h130e100c;
	16'h807 : data <= 32'h93001000;
	16'h808 : data <= 32'h13010000;
	16'h809 : data <= 32'h63e42000;
	16'h80a : data <= 32'h6316c001;
	16'h80b : data <= 32'h6304c001;
	16'h80c : data <= 32'h6f505022;
	16'h80d : data <= 32'he3ec20fe;
	16'h80e : data <= 32'h130e200c;
	16'h80f : data <= 32'h9300f0ff;
	16'h810 : data <= 32'h1301e0ff;
	16'h811 : data <= 32'h63e42000;
	16'h812 : data <= 32'h6316c001;
	16'h813 : data <= 32'h6304c001;
	16'h814 : data <= 32'h6f505020;
	16'h815 : data <= 32'he3ec20fe;
	16'h816 : data <= 32'h130e300c;
	16'h817 : data <= 32'h9300f0ff;
	16'h818 : data <= 32'h13010000;
	16'h819 : data <= 32'h63e42000;
	16'h81a : data <= 32'h6316c001;
	16'h81b : data <= 32'h6304c001;
	16'h81c : data <= 32'h6f50501e;
	16'h81d : data <= 32'he3ec20fe;
	16'h81e : data <= 32'h130e400c;
	16'h81f : data <= 32'hb7000080;
	16'h820 : data <= 32'h37010080;
	16'h821 : data <= 32'h1301f1ff;
	16'h822 : data <= 32'h63e42000;
	16'h823 : data <= 32'h6316c001;
	16'h824 : data <= 32'h6304c001;
	16'h825 : data <= 32'h6f50101c;
	16'h826 : data <= 32'he3ec20fe;
	16'h827 : data <= 32'h130e500c;
	16'h828 : data <= 32'h13020000;
	16'h829 : data <= 32'hb70000f0;
	16'h82a : data <= 32'h370100f0;
	16'h82b : data <= 32'h1301f1ff;
	16'h82c : data <= 32'h63f42000;
	16'h82d : data <= 32'h6f50101a;
	16'h82e : data <= 32'h13021200;
	16'h82f : data <= 32'h93022000;
	16'h830 : data <= 32'he31252fe;
	16'h831 : data <= 32'h130e600c;
	16'h832 : data <= 32'h13020000;
	16'h833 : data <= 32'hb70000f0;
	16'h834 : data <= 32'h370100f0;
	16'h835 : data <= 32'h1301f1ff;
	16'h836 : data <= 32'h13000000;
	16'h837 : data <= 32'h63f42000;
	16'h838 : data <= 32'h6f505017;
	16'h839 : data <= 32'h13021200;
	16'h83a : data <= 32'h93022000;
	16'h83b : data <= 32'he31052fe;
	16'h83c : data <= 32'h130e700c;
	16'h83d : data <= 32'h13020000;
	16'h83e : data <= 32'hb70000f0;
	16'h83f : data <= 32'h370100f0;
	16'h840 : data <= 32'h1301f1ff;
	16'h841 : data <= 32'h13000000;
	16'h842 : data <= 32'h13000000;
	16'h843 : data <= 32'h63f42000;
	16'h844 : data <= 32'h6f505014;
	16'h845 : data <= 32'h13021200;
	16'h846 : data <= 32'h93022000;
	16'h847 : data <= 32'he31e52fc;
	16'h848 : data <= 32'h130e800c;
	16'h849 : data <= 32'h13020000;
	16'h84a : data <= 32'hb70000f0;
	16'h84b : data <= 32'h13000000;
	16'h84c : data <= 32'h370100f0;
	16'h84d : data <= 32'h1301f1ff;
	16'h84e : data <= 32'h63f42000;
	16'h84f : data <= 32'h6f509011;
	16'h850 : data <= 32'h13021200;
	16'h851 : data <= 32'h93022000;
	16'h852 : data <= 32'he31052fe;
	16'h853 : data <= 32'h130e900c;
	16'h854 : data <= 32'h13020000;
	16'h855 : data <= 32'hb70000f0;
	16'h856 : data <= 32'h13000000;
	16'h857 : data <= 32'h370100f0;
	16'h858 : data <= 32'h1301f1ff;
	16'h859 : data <= 32'h13000000;
	16'h85a : data <= 32'h63f42000;
	16'h85b : data <= 32'h6f50900e;
	16'h85c : data <= 32'h13021200;
	16'h85d : data <= 32'h93022000;
	16'h85e : data <= 32'he31e52fc;
	16'h85f : data <= 32'h130ea00c;
	16'h860 : data <= 32'h13020000;
	16'h861 : data <= 32'hb70000f0;
	16'h862 : data <= 32'h13000000;
	16'h863 : data <= 32'h13000000;
	16'h864 : data <= 32'h370100f0;
	16'h865 : data <= 32'h1301f1ff;
	16'h866 : data <= 32'h63f42000;
	16'h867 : data <= 32'h6f50900b;
	16'h868 : data <= 32'h13021200;
	16'h869 : data <= 32'h93022000;
	16'h86a : data <= 32'he31e52fc;
	16'h86b : data <= 32'h130eb00c;
	16'h86c : data <= 32'h13020000;
	16'h86d : data <= 32'hb70000f0;
	16'h86e : data <= 32'h370100f0;
	16'h86f : data <= 32'h1301f1ff;
	16'h870 : data <= 32'h63f42000;
	16'h871 : data <= 32'h6f501009;
	16'h872 : data <= 32'h13021200;
	16'h873 : data <= 32'h93022000;
	16'h874 : data <= 32'he31252fe;
	16'h875 : data <= 32'h130ec00c;
	16'h876 : data <= 32'h13020000;
	16'h877 : data <= 32'hb70000f0;
	16'h878 : data <= 32'h370100f0;
	16'h879 : data <= 32'h1301f1ff;
	16'h87a : data <= 32'h13000000;
	16'h87b : data <= 32'h63f42000;
	16'h87c : data <= 32'h6f505006;
	16'h87d : data <= 32'h13021200;
	16'h87e : data <= 32'h93022000;
	16'h87f : data <= 32'he31052fe;
	16'h880 : data <= 32'h130ed00c;
	16'h881 : data <= 32'h13020000;
	16'h882 : data <= 32'hb70000f0;
	16'h883 : data <= 32'h370100f0;
	16'h884 : data <= 32'h1301f1ff;
	16'h885 : data <= 32'h13000000;
	16'h886 : data <= 32'h13000000;
	16'h887 : data <= 32'h63f42000;
	16'h888 : data <= 32'h6f505003;
	16'h889 : data <= 32'h13021200;
	16'h88a : data <= 32'h93022000;
	16'h88b : data <= 32'he31e52fc;
	16'h88c : data <= 32'h130ee00c;
	16'h88d : data <= 32'h13020000;
	16'h88e : data <= 32'hb70000f0;
	16'h88f : data <= 32'h13000000;
	16'h890 : data <= 32'h370100f0;
	16'h891 : data <= 32'h1301f1ff;
	16'h892 : data <= 32'h63f42000;
	16'h893 : data <= 32'h6f509000;
	16'h894 : data <= 32'h13021200;
	16'h895 : data <= 32'h93022000;
	16'h896 : data <= 32'he31052fe;
	16'h897 : data <= 32'h130ef00c;
	16'h898 : data <= 32'h13020000;
	16'h899 : data <= 32'hb70000f0;
	16'h89a : data <= 32'h13000000;
	16'h89b : data <= 32'h370100f0;
	16'h89c : data <= 32'h1301f1ff;
	16'h89d : data <= 32'h13000000;
	16'h89e : data <= 32'h63f42000;
	16'h89f : data <= 32'h6f50807d;
	16'h8a0 : data <= 32'h13021200;
	16'h8a1 : data <= 32'h93022000;
	16'h8a2 : data <= 32'he31e52fc;
	16'h8a3 : data <= 32'h130e000d;
	16'h8a4 : data <= 32'h13020000;
	16'h8a5 : data <= 32'hb70000f0;
	16'h8a6 : data <= 32'h13000000;
	16'h8a7 : data <= 32'h13000000;
	16'h8a8 : data <= 32'h370100f0;
	16'h8a9 : data <= 32'h1301f1ff;
	16'h8aa : data <= 32'h63f42000;
	16'h8ab : data <= 32'h6f50807a;
	16'h8ac : data <= 32'h13021200;
	16'h8ad : data <= 32'h93022000;
	16'h8ae : data <= 32'he31e52fc;
	16'h8af : data <= 32'h93001000;
	16'h8b0 : data <= 32'h636a1000;
	16'h8b1 : data <= 32'h93801000;
	16'h8b2 : data <= 32'h93801000;
	16'h8b3 : data <= 32'h93801000;
	16'h8b4 : data <= 32'h93801000;
	16'h8b5 : data <= 32'h93801000;
	16'h8b6 : data <= 32'h93801000;
	16'h8b7 : data <= 32'h930e3000;
	16'h8b8 : data <= 32'h130e100d;
	16'h8b9 : data <= 32'h6384d001;
	16'h8ba : data <= 32'h6f50c076;
	16'h8bb : data <= 32'h130e200d;
	16'h8bc : data <= 32'h93000000;
	16'h8bd : data <= 32'h13011000;
	16'h8be : data <= 32'h63982000;
	16'h8bf : data <= 32'h6304c001;
	16'h8c0 : data <= 32'h6f504075;
	16'h8c1 : data <= 32'h6318c001;
	16'h8c2 : data <= 32'he39e20fe;
	16'h8c3 : data <= 32'h6304c001;
	16'h8c4 : data <= 32'h6f504074;
	16'h8c5 : data <= 32'h130e300d;
	16'h8c6 : data <= 32'h93001000;
	16'h8c7 : data <= 32'h13010000;
	16'h8c8 : data <= 32'h63982000;
	16'h8c9 : data <= 32'h6304c001;
	16'h8ca : data <= 32'h6f50c072;
	16'h8cb : data <= 32'h6318c001;
	16'h8cc : data <= 32'he39e20fe;
	16'h8cd : data <= 32'h6304c001;
	16'h8ce : data <= 32'h6f50c071;
	16'h8cf : data <= 32'h130e400d;
	16'h8d0 : data <= 32'h9300f0ff;
	16'h8d1 : data <= 32'h13011000;
	16'h8d2 : data <= 32'h63982000;
	16'h8d3 : data <= 32'h6304c001;
	16'h8d4 : data <= 32'h6f504070;
	16'h8d5 : data <= 32'h6318c001;
	16'h8d6 : data <= 32'he39e20fe;
	16'h8d7 : data <= 32'h6304c001;
	16'h8d8 : data <= 32'h6f50406f;
	16'h8d9 : data <= 32'h130e500d;
	16'h8da : data <= 32'h93001000;
	16'h8db : data <= 32'h1301f0ff;
	16'h8dc : data <= 32'h63982000;
	16'h8dd : data <= 32'h6304c001;
	16'h8de : data <= 32'h6f50c06d;
	16'h8df : data <= 32'h6318c001;
	16'h8e0 : data <= 32'he39e20fe;
	16'h8e1 : data <= 32'h6304c001;
	16'h8e2 : data <= 32'h6f50c06c;
	16'h8e3 : data <= 32'h130e600d;
	16'h8e4 : data <= 32'h93000000;
	16'h8e5 : data <= 32'h13010000;
	16'h8e6 : data <= 32'h63942000;
	16'h8e7 : data <= 32'h6316c001;
	16'h8e8 : data <= 32'h6304c001;
	16'h8e9 : data <= 32'h6f50006b;
	16'h8ea : data <= 32'he39c20fe;
	16'h8eb : data <= 32'h130e700d;
	16'h8ec : data <= 32'h93001000;
	16'h8ed : data <= 32'h13011000;
	16'h8ee : data <= 32'h63942000;
	16'h8ef : data <= 32'h6316c001;
	16'h8f0 : data <= 32'h6304c001;
	16'h8f1 : data <= 32'h6f500069;
	16'h8f2 : data <= 32'he39c20fe;
	16'h8f3 : data <= 32'h130e800d;
	16'h8f4 : data <= 32'h9300f0ff;
	16'h8f5 : data <= 32'h1301f0ff;
	16'h8f6 : data <= 32'h63942000;
	16'h8f7 : data <= 32'h6316c001;
	16'h8f8 : data <= 32'h6304c001;
	16'h8f9 : data <= 32'h6f500067;
	16'h8fa : data <= 32'he39c20fe;
	16'h8fb : data <= 32'h130e900d;
	16'h8fc : data <= 32'h13020000;
	16'h8fd : data <= 32'h93000000;
	16'h8fe : data <= 32'h13010000;
	16'h8ff : data <= 32'h63842000;
	16'h900 : data <= 32'h6f504065;
	16'h901 : data <= 32'h13021200;
	16'h902 : data <= 32'h93022000;
	16'h903 : data <= 32'he31452fe;
	16'h904 : data <= 32'h130ea00d;
	16'h905 : data <= 32'h13020000;
	16'h906 : data <= 32'h93000000;
	16'h907 : data <= 32'h13010000;
	16'h908 : data <= 32'h13000000;
	16'h909 : data <= 32'h63842000;
	16'h90a : data <= 32'h6f50c062;
	16'h90b : data <= 32'h13021200;
	16'h90c : data <= 32'h93022000;
	16'h90d : data <= 32'he31252fe;
	16'h90e : data <= 32'h130eb00d;
	16'h90f : data <= 32'h13020000;
	16'h910 : data <= 32'h93000000;
	16'h911 : data <= 32'h13010000;
	16'h912 : data <= 32'h13000000;
	16'h913 : data <= 32'h13000000;
	16'h914 : data <= 32'h63842000;
	16'h915 : data <= 32'h6f500060;
	16'h916 : data <= 32'h13021200;
	16'h917 : data <= 32'h93022000;
	16'h918 : data <= 32'he31052fe;
	16'h919 : data <= 32'h130ec00d;
	16'h91a : data <= 32'h13020000;
	16'h91b : data <= 32'h93000000;
	16'h91c : data <= 32'h13000000;
	16'h91d : data <= 32'h13010000;
	16'h91e : data <= 32'h63842000;
	16'h91f : data <= 32'h6f50805d;
	16'h920 : data <= 32'h13021200;
	16'h921 : data <= 32'h93022000;
	16'h922 : data <= 32'he31252fe;
	16'h923 : data <= 32'h130ed00d;
	16'h924 : data <= 32'h13020000;
	16'h925 : data <= 32'h93000000;
	16'h926 : data <= 32'h13000000;
	16'h927 : data <= 32'h13010000;
	16'h928 : data <= 32'h13000000;
	16'h929 : data <= 32'h63842000;
	16'h92a : data <= 32'h6f50c05a;
	16'h92b : data <= 32'h13021200;
	16'h92c : data <= 32'h93022000;
	16'h92d : data <= 32'he31052fe;
	16'h92e : data <= 32'h130ee00d;
	16'h92f : data <= 32'h13020000;
	16'h930 : data <= 32'h93000000;
	16'h931 : data <= 32'h13000000;
	16'h932 : data <= 32'h13000000;
	16'h933 : data <= 32'h13010000;
	16'h934 : data <= 32'h63842000;
	16'h935 : data <= 32'h6f500058;
	16'h936 : data <= 32'h13021200;
	16'h937 : data <= 32'h93022000;
	16'h938 : data <= 32'he31052fe;
	16'h939 : data <= 32'h130ef00d;
	16'h93a : data <= 32'h13020000;
	16'h93b : data <= 32'h93000000;
	16'h93c : data <= 32'h13010000;
	16'h93d : data <= 32'h63842000;
	16'h93e : data <= 32'h6f50c055;
	16'h93f : data <= 32'h13021200;
	16'h940 : data <= 32'h93022000;
	16'h941 : data <= 32'he31452fe;
	16'h942 : data <= 32'h130e000e;
	16'h943 : data <= 32'h13020000;
	16'h944 : data <= 32'h93000000;
	16'h945 : data <= 32'h13010000;
	16'h946 : data <= 32'h13000000;
	16'h947 : data <= 32'h63842000;
	16'h948 : data <= 32'h6f504053;
	16'h949 : data <= 32'h13021200;
	16'h94a : data <= 32'h93022000;
	16'h94b : data <= 32'he31252fe;
	16'h94c : data <= 32'h130e100e;
	16'h94d : data <= 32'h13020000;
	16'h94e : data <= 32'h93000000;
	16'h94f : data <= 32'h13010000;
	16'h950 : data <= 32'h13000000;
	16'h951 : data <= 32'h13000000;
	16'h952 : data <= 32'h63842000;
	16'h953 : data <= 32'h6f508050;
	16'h954 : data <= 32'h13021200;
	16'h955 : data <= 32'h93022000;
	16'h956 : data <= 32'he31052fe;
	16'h957 : data <= 32'h130e200e;
	16'h958 : data <= 32'h13020000;
	16'h959 : data <= 32'h93000000;
	16'h95a : data <= 32'h13000000;
	16'h95b : data <= 32'h13010000;
	16'h95c : data <= 32'h63842000;
	16'h95d : data <= 32'h6f50004e;
	16'h95e : data <= 32'h13021200;
	16'h95f : data <= 32'h93022000;
	16'h960 : data <= 32'he31252fe;
	16'h961 : data <= 32'h130e300e;
	16'h962 : data <= 32'h13020000;
	16'h963 : data <= 32'h93000000;
	16'h964 : data <= 32'h13000000;
	16'h965 : data <= 32'h13010000;
	16'h966 : data <= 32'h13000000;
	16'h967 : data <= 32'h63842000;
	16'h968 : data <= 32'h6f50404b;
	16'h969 : data <= 32'h13021200;
	16'h96a : data <= 32'h93022000;
	16'h96b : data <= 32'he31052fe;
	16'h96c : data <= 32'h130e400e;
	16'h96d : data <= 32'h13020000;
	16'h96e : data <= 32'h93000000;
	16'h96f : data <= 32'h13000000;
	16'h970 : data <= 32'h13000000;
	16'h971 : data <= 32'h13010000;
	16'h972 : data <= 32'h63842000;
	16'h973 : data <= 32'h6f508048;
	16'h974 : data <= 32'h13021200;
	16'h975 : data <= 32'h93022000;
	16'h976 : data <= 32'he31052fe;
	16'h977 : data <= 32'h93001000;
	16'h978 : data <= 32'h639a0000;
	16'h979 : data <= 32'h93801000;
	16'h97a : data <= 32'h93801000;
	16'h97b : data <= 32'h93801000;
	16'h97c : data <= 32'h93801000;
	16'h97d : data <= 32'h93801000;
	16'h97e : data <= 32'h93801000;
	16'h97f : data <= 32'h930e3000;
	16'h980 : data <= 32'h130e500e;
	16'h981 : data <= 32'h6384d001;
	16'h982 : data <= 32'h6f50c044;
	16'h983 : data <= 32'h73100034;
	16'h984 : data <= 32'h9360000f;
	16'h985 : data <= 32'h1361f000;
	16'h986 : data <= 32'h93611000;
	16'h987 : data <= 32'h1362f00f;
	16'h988 : data <= 32'hf3a10034;
	16'h989 : data <= 32'h63123002;
	16'h98a : data <= 32'h93611000;
	16'h98b : data <= 32'hf3210034;
	16'h98c : data <= 32'h639c1100;
	16'h98d : data <= 32'hf3210134;
	16'h98e : data <= 32'h63981100;
	16'h98f : data <= 32'h0f00f00f;
	16'h990 : data <= 32'h130e1000;
	16'h991 : data <= 32'h6f500043;
	16'h992 : data <= 32'h0f00f00f;
	16'h993 : data <= 32'h63000e00;
	16'h994 : data <= 32'h131e1e00;
	16'h995 : data <= 32'h136e1e00;
	16'h996 : data <= 32'h6f50c041;
	16'h997 : data <= 32'h9306f006;
	16'h998 : data <= 32'h17050000;
	16'h999 : data <= 32'h13058507;
	16'h99a : data <= 32'h97050000;
	16'h99b : data <= 32'h93850502;
	16'h99c : data <= 32'h17060000;
	16'h99d : data <= 32'h13060605;
	16'h99e : data <= 32'h03250500;
	16'h99f : data <= 32'h13000000;
	16'h9a0 : data <= 32'h23a0a500;
	16'h9a1 : data <= 32'h0f100000;
	16'h9a2 : data <= 32'h9386e60d;
	16'h9a3 : data <= 32'h13000000;
	16'h9a4 : data <= 32'h930ec01b;
	16'h9a5 : data <= 32'h130e600e;
	16'h9a6 : data <= 32'h6384d601;
	16'h9a7 : data <= 32'h6f50803b;
	16'h9a8 : data <= 32'h13074006;
	16'h9a9 : data <= 32'h1307f7ff;
	16'h9aa : data <= 32'he31e07fe;
	16'h9ab : data <= 32'h2320a600;
	16'h9ac : data <= 32'h0f100000;
	16'h9ad : data <= 32'h13000000;
	16'h9ae : data <= 32'h13000000;
	16'h9af : data <= 32'h13000000;
	16'h9b0 : data <= 32'h9386b622;
	16'h9b1 : data <= 32'h13000000;
	16'h9b2 : data <= 32'h930e9030;
	16'h9b3 : data <= 32'h130e700e;
	16'h9b4 : data <= 32'h6384d601;
	16'h9b5 : data <= 32'h6f500038;
	16'h9b6 : data <= 32'h9386d614;
	16'h9b7 : data <= 32'h130e800e;
	16'h9b8 : data <= 32'h6f008000;
	16'h9b9 : data <= 32'h6f500037;
	16'h9ba : data <= 32'h93001000;
	16'h9bb : data <= 32'h6f004001;
	16'h9bc : data <= 32'h93801000;
	16'h9bd : data <= 32'h93801000;
	16'h9be : data <= 32'h93801000;
	16'h9bf : data <= 32'h93801000;
	16'h9c0 : data <= 32'h93801000;
	16'h9c1 : data <= 32'h93801000;
	16'h9c2 : data <= 32'h930e3000;
	16'h9c3 : data <= 32'h130e900e;
	16'h9c4 : data <= 32'h6384d001;
	16'h9c5 : data <= 32'h6f500034;
	16'h9c6 : data <= 32'h130ea00e;
	16'h9c7 : data <= 32'h93000000;
	16'h9c8 : data <= 32'hef000001;
	16'h9c9 : data <= 32'h13000000;
	16'h9ca : data <= 32'h13000000;
	16'h9cb : data <= 32'h6f508032;
	16'h9cc : data <= 32'h17010000;
	16'h9cd : data <= 32'h130101ff;
	16'h9ce : data <= 32'h13014100;
	16'h9cf : data <= 32'h63041100;
	16'h9d0 : data <= 32'h6f504031;
	16'h9d1 : data <= 32'h13011000;
	16'h9d2 : data <= 32'hef004001;
	16'h9d3 : data <= 32'h13011100;
	16'h9d4 : data <= 32'h13011100;
	16'h9d5 : data <= 32'h13011100;
	16'h9d6 : data <= 32'h13011100;
	16'h9d7 : data <= 32'h13011100;
	16'h9d8 : data <= 32'h13011100;
	16'h9d9 : data <= 32'h930e3000;
	16'h9da : data <= 32'h130eb00e;
	16'h9db : data <= 32'h6304d101;
	16'h9dc : data <= 32'h6f50402e;
	16'h9dd : data <= 32'h130ec00e;
	16'h9de : data <= 32'h930f0000;
	16'h9df : data <= 32'h17010000;
	16'h9e0 : data <= 32'h13018101;
	16'h9e1 : data <= 32'he7090100;
	16'h9e2 : data <= 32'h13000000;
	16'h9e3 : data <= 32'h13000000;
	16'h9e4 : data <= 32'h6f50402c;
	16'h9e5 : data <= 32'h97000000;
	16'h9e6 : data <= 32'h938000ff;
	16'h9e7 : data <= 32'h93804000;
	16'h9e8 : data <= 32'h63843001;
	16'h9e9 : data <= 32'h6f50002b;
	16'h9ea : data <= 32'h130ed00e;
	16'h9eb : data <= 32'h930f0000;
	16'h9ec : data <= 32'h97010000;
	16'h9ed : data <= 32'h93814101;
	16'h9ee : data <= 32'h67800100;
	16'h9ef : data <= 32'h13000000;
	16'h9f0 : data <= 32'h6f504029;
	16'h9f1 : data <= 32'h63840f00;
	16'h9f2 : data <= 32'h6f50c028;
	16'h9f3 : data <= 32'h130ee00e;
	16'h9f4 : data <= 32'h13020000;
	16'h9f5 : data <= 32'h17030000;
	16'h9f6 : data <= 32'h13034301;
	16'h9f7 : data <= 32'he7090300;
	16'h9f8 : data <= 32'h6304c001;
	16'h9f9 : data <= 32'h6f500027;
	16'h9fa : data <= 32'h13021200;
	16'h9fb : data <= 32'h93022000;
	16'h9fc : data <= 32'he31252fe;
	16'h9fd : data <= 32'h130ef00e;
	16'h9fe : data <= 32'h13020000;
	16'h9ff : data <= 32'h17030000;
	16'ha00 : data <= 32'h13038301;
	16'ha01 : data <= 32'h13000000;
	16'ha02 : data <= 32'he7090300;
	16'ha03 : data <= 32'h6304c001;
	16'ha04 : data <= 32'h6f504024;
	16'ha05 : data <= 32'h13021200;
	16'ha06 : data <= 32'h93022000;
	16'ha07 : data <= 32'he31052fe;
	16'ha08 : data <= 32'h130e000f;
	16'ha09 : data <= 32'h13020000;
	16'ha0a : data <= 32'h17030000;
	16'ha0b : data <= 32'h1303c301;
	16'ha0c : data <= 32'h13000000;
	16'ha0d : data <= 32'h13000000;
	16'ha0e : data <= 32'he7090300;
	16'ha0f : data <= 32'h6304c001;
	16'ha10 : data <= 32'h6f504021;
	16'ha11 : data <= 32'h13021200;
	16'ha12 : data <= 32'h93022000;
	16'ha13 : data <= 32'he31e52fc;
	16'ha14 : data <= 32'h93001000;
	16'ha15 : data <= 32'h17010000;
	16'ha16 : data <= 32'h1301c101;
	16'ha17 : data <= 32'he709c1ff;
	16'ha18 : data <= 32'h93801000;
	16'ha19 : data <= 32'h93801000;
	16'ha1a : data <= 32'h93801000;
	16'ha1b : data <= 32'h93801000;
	16'ha1c : data <= 32'h93801000;
	16'ha1d : data <= 32'h93801000;
	16'ha1e : data <= 32'h930e4000;
	16'ha1f : data <= 32'h130e100f;
	16'ha20 : data <= 32'h6384d001;
	16'ha21 : data <= 32'h6f50001d;
	16'ha22 : data <= 32'h97500000;
	16'ha23 : data <= 32'h93808077;
	16'ha24 : data <= 32'h83810000;
	16'ha25 : data <= 32'h930ef0ff;
	16'ha26 : data <= 32'h130e200f;
	16'ha27 : data <= 32'h6384d101;
	16'ha28 : data <= 32'h6f50401b;
	16'ha29 : data <= 32'h97500000;
	16'ha2a : data <= 32'h9380c075;
	16'ha2b : data <= 32'h83811000;
	16'ha2c : data <= 32'h930e0000;
	16'ha2d : data <= 32'h130e300f;
	16'ha2e : data <= 32'h6384d101;
	16'ha2f : data <= 32'h6f508019;
	16'ha30 : data <= 32'h97500000;
	16'ha31 : data <= 32'h93800074;
	16'ha32 : data <= 32'h83812000;
	16'ha33 : data <= 32'h930e00ff;
	16'ha34 : data <= 32'h130e400f;
	16'ha35 : data <= 32'h6384d101;
	16'ha36 : data <= 32'h6f50c017;
	16'ha37 : data <= 32'h97500000;
	16'ha38 : data <= 32'h93804072;
	16'ha39 : data <= 32'h83813000;
	16'ha3a : data <= 32'h930ef000;
	16'ha3b : data <= 32'h130e500f;
	16'ha3c : data <= 32'h6384d101;
	16'ha3d : data <= 32'h6f500016;
	16'ha3e : data <= 32'h97500000;
	16'ha3f : data <= 32'h9380b070;
	16'ha40 : data <= 32'h8381d0ff;
	16'ha41 : data <= 32'h930ef0ff;
	16'ha42 : data <= 32'h130e600f;
	16'ha43 : data <= 32'h6384d101;
	16'ha44 : data <= 32'h6f504014;
	16'ha45 : data <= 32'h97500000;
	16'ha46 : data <= 32'h9380f06e;
	16'ha47 : data <= 32'h8381e0ff;
	16'ha48 : data <= 32'h930e0000;
	16'ha49 : data <= 32'h130e700f;
	16'ha4a : data <= 32'h6384d101;
	16'ha4b : data <= 32'h6f508012;
	16'ha4c : data <= 32'h97500000;
	16'ha4d : data <= 32'h9380306d;
	16'ha4e : data <= 32'h8381f0ff;
	16'ha4f : data <= 32'h930e00ff;
	16'ha50 : data <= 32'h130e800f;
	16'ha51 : data <= 32'h6384d101;
	16'ha52 : data <= 32'h6f50c010;
	16'ha53 : data <= 32'h97500000;
	16'ha54 : data <= 32'h9380706b;
	16'ha55 : data <= 32'h83810000;
	16'ha56 : data <= 32'h930ef000;
	16'ha57 : data <= 32'h130e900f;
	16'ha58 : data <= 32'h6384d101;
	16'ha59 : data <= 32'h6f50000f;
	16'ha5a : data <= 32'h97500000;
	16'ha5b : data <= 32'h93808069;
	16'ha5c : data <= 32'h938000fe;
	16'ha5d : data <= 32'h83810002;
	16'ha5e : data <= 32'h930ef0ff;
	16'ha5f : data <= 32'h130ea00f;
	16'ha60 : data <= 32'h6384d101;
	16'ha61 : data <= 32'h6f50000d;
	16'ha62 : data <= 32'h97500000;
	16'ha63 : data <= 32'h93808067;
	16'ha64 : data <= 32'h9380a0ff;
	16'ha65 : data <= 32'h83817000;
	16'ha66 : data <= 32'h930e0000;
	16'ha67 : data <= 32'h130eb00f;
	16'ha68 : data <= 32'h6384d101;
	16'ha69 : data <= 32'h6f50000b;
	16'ha6a : data <= 32'h130ec00f;
	16'ha6b : data <= 32'h13020000;
	16'ha6c : data <= 32'h97500000;
	16'ha6d : data <= 32'h93801065;
	16'ha6e : data <= 32'h83811000;
	16'ha6f : data <= 32'h13830100;
	16'ha70 : data <= 32'h930e00ff;
	16'ha71 : data <= 32'h6304d301;
	16'ha72 : data <= 32'h6f50c008;
	16'ha73 : data <= 32'h13021200;
	16'ha74 : data <= 32'h93022000;
	16'ha75 : data <= 32'he31e52fc;
	16'ha76 : data <= 32'h130ed00f;
	16'ha77 : data <= 32'h13020000;
	16'ha78 : data <= 32'h97500000;
	16'ha79 : data <= 32'h93802062;
	16'ha7a : data <= 32'h83811000;
	16'ha7b : data <= 32'h13000000;
	16'ha7c : data <= 32'h13830100;
	16'ha7d : data <= 32'h930ef000;
	16'ha7e : data <= 32'h6304d301;
	16'ha7f : data <= 32'h6f508005;
	16'ha80 : data <= 32'h13021200;
	16'ha81 : data <= 32'h93022000;
	16'ha82 : data <= 32'he31c52fc;
	16'ha83 : data <= 32'h130ee00f;
	16'ha84 : data <= 32'h13020000;
	16'ha85 : data <= 32'h97500000;
	16'ha86 : data <= 32'h9380c05e;
	16'ha87 : data <= 32'h83811000;
	16'ha88 : data <= 32'h13000000;
	16'ha89 : data <= 32'h13000000;
	16'ha8a : data <= 32'h13830100;
	16'ha8b : data <= 32'h930e0000;
	16'ha8c : data <= 32'h6304d301;
	16'ha8d : data <= 32'h6f500002;
	16'ha8e : data <= 32'h13021200;
	16'ha8f : data <= 32'h93022000;
	16'ha90 : data <= 32'he31a52fc;
	16'ha91 : data <= 32'h130ef00f;
	16'ha92 : data <= 32'h13020000;
	16'ha93 : data <= 32'h97500000;
	16'ha94 : data <= 32'h9380505b;
	16'ha95 : data <= 32'h83811000;
	16'ha96 : data <= 32'h930e00ff;
	16'ha97 : data <= 32'h6384d101;
	16'ha98 : data <= 32'h6f40507f;
	16'ha99 : data <= 32'h13021200;
	16'ha9a : data <= 32'h93022000;
	16'ha9b : data <= 32'he31052fe;
	16'ha9c : data <= 32'h130e0010;
	16'ha9d : data <= 32'h13020000;
	16'ha9e : data <= 32'h97500000;
	16'ha9f : data <= 32'h9380a058;
	16'haa0 : data <= 32'h13000000;
	16'haa1 : data <= 32'h83811000;
	16'haa2 : data <= 32'h930ef000;
	16'haa3 : data <= 32'h6384d101;
	16'haa4 : data <= 32'h6f40507c;
	16'haa5 : data <= 32'h13021200;
	16'haa6 : data <= 32'h93022000;
	16'haa7 : data <= 32'he31e52fc;
	16'haa8 : data <= 32'h130e1010;
	16'haa9 : data <= 32'h13020000;
	16'haaa : data <= 32'h97500000;
	16'haab : data <= 32'h93808055;
	16'haac : data <= 32'h13000000;
	16'haad : data <= 32'h13000000;
	16'haae : data <= 32'h83811000;
	16'haaf : data <= 32'h930e0000;
	16'hab0 : data <= 32'h6384d101;
	16'hab1 : data <= 32'h6f401079;
	16'hab2 : data <= 32'h13021200;
	16'hab3 : data <= 32'h93022000;
	16'hab4 : data <= 32'he31c52fc;
	16'hab5 : data <= 32'h97510000;
	16'hab6 : data <= 32'h9381c152;
	16'hab7 : data <= 32'h03810100;
	16'hab8 : data <= 32'h13012000;
	16'hab9 : data <= 32'h930e2000;
	16'haba : data <= 32'h130e2010;
	16'habb : data <= 32'h6304d101;
	16'habc : data <= 32'h6f405076;
	16'habd : data <= 32'h97510000;
	16'habe : data <= 32'h9381c150;
	16'habf : data <= 32'h03810100;
	16'hac0 : data <= 32'h13000000;
	16'hac1 : data <= 32'h13012000;
	16'hac2 : data <= 32'h930e2000;
	16'hac3 : data <= 32'h130e3010;
	16'hac4 : data <= 32'h6304d101;
	16'hac5 : data <= 32'h6f401074;
	16'hac6 : data <= 32'h97500000;
	16'hac7 : data <= 32'h9380c04e;
	16'hac8 : data <= 32'h83c10000;
	16'hac9 : data <= 32'h930ef00f;
	16'haca : data <= 32'h130e4010;
	16'hacb : data <= 32'h6384d101;
	16'hacc : data <= 32'h6f405072;
	16'hacd : data <= 32'h97500000;
	16'hace : data <= 32'h9380004d;
	16'hacf : data <= 32'h83c11000;
	16'had0 : data <= 32'h930e0000;
	16'had1 : data <= 32'h130e5010;
	16'had2 : data <= 32'h6384d101;
	16'had3 : data <= 32'h6f409070;
	16'had4 : data <= 32'h97500000;
	16'had5 : data <= 32'h9380404b;
	16'had6 : data <= 32'h83c12000;
	16'had7 : data <= 32'h930e000f;
	16'had8 : data <= 32'h130e6010;
	16'had9 : data <= 32'h6384d101;
	16'hada : data <= 32'h6f40d06e;
	16'hadb : data <= 32'h97500000;
	16'hadc : data <= 32'h93808049;
	16'hadd : data <= 32'h83c13000;
	16'hade : data <= 32'h930ef000;
	16'hadf : data <= 32'h130e7010;
	16'hae0 : data <= 32'h6384d101;
	16'hae1 : data <= 32'h6f40106d;
	16'hae2 : data <= 32'h97500000;
	16'hae3 : data <= 32'h9380f047;
	16'hae4 : data <= 32'h83c1d0ff;
	16'hae5 : data <= 32'h930ef00f;
	16'hae6 : data <= 32'h130e8010;
	16'hae7 : data <= 32'h6384d101;
	16'hae8 : data <= 32'h6f40506b;
	16'hae9 : data <= 32'h97500000;
	16'haea : data <= 32'h93803046;
	16'haeb : data <= 32'h83c1e0ff;
	16'haec : data <= 32'h930e0000;
	16'haed : data <= 32'h130e9010;
	16'haee : data <= 32'h6384d101;
	16'haef : data <= 32'h6f409069;
	16'haf0 : data <= 32'h97500000;
	16'haf1 : data <= 32'h93807044;
	16'haf2 : data <= 32'h83c1f0ff;
	16'haf3 : data <= 32'h930e000f;
	16'haf4 : data <= 32'h130ea010;
	16'haf5 : data <= 32'h6384d101;
	16'haf6 : data <= 32'h6f40d067;
	16'haf7 : data <= 32'h97500000;
	16'haf8 : data <= 32'h9380b042;
	16'haf9 : data <= 32'h83c10000;
	16'hafa : data <= 32'h930ef000;
	16'hafb : data <= 32'h130eb010;
	16'hafc : data <= 32'h6384d101;
	16'hafd : data <= 32'h6f401066;
	16'hafe : data <= 32'h97500000;
	16'haff : data <= 32'h9380c040;
	16'hb00 : data <= 32'h938000fe;
	16'hb01 : data <= 32'h83c10002;
	16'hb02 : data <= 32'h930ef00f;
	16'hb03 : data <= 32'h130ec010;
	16'hb04 : data <= 32'h6384d101;
	16'hb05 : data <= 32'h6f401064;
	16'hb06 : data <= 32'h97500000;
	16'hb07 : data <= 32'h9380c03e;
	16'hb08 : data <= 32'h9380a0ff;
	16'hb09 : data <= 32'h83c17000;
	16'hb0a : data <= 32'h930e0000;
	16'hb0b : data <= 32'h130ed010;
	16'hb0c : data <= 32'h6384d101;
	16'hb0d : data <= 32'h6f401062;
	16'hb0e : data <= 32'h130ee010;
	16'hb0f : data <= 32'h13020000;
	16'hb10 : data <= 32'h97500000;
	16'hb11 : data <= 32'h9380503c;
	16'hb12 : data <= 32'h83c11000;
	16'hb13 : data <= 32'h13830100;
	16'hb14 : data <= 32'h930e000f;
	16'hb15 : data <= 32'h6304d301;
	16'hb16 : data <= 32'h6f40d05f;
	16'hb17 : data <= 32'h13021200;
	16'hb18 : data <= 32'h93022000;
	16'hb19 : data <= 32'he31e52fc;
	16'hb1a : data <= 32'h130ef010;
	16'hb1b : data <= 32'h13020000;
	16'hb1c : data <= 32'h97500000;
	16'hb1d : data <= 32'h93806039;
	16'hb1e : data <= 32'h83c11000;
	16'hb1f : data <= 32'h13000000;
	16'hb20 : data <= 32'h13830100;
	16'hb21 : data <= 32'h930ef000;
	16'hb22 : data <= 32'h6304d301;
	16'hb23 : data <= 32'h6f40905c;
	16'hb24 : data <= 32'h13021200;
	16'hb25 : data <= 32'h93022000;
	16'hb26 : data <= 32'he31c52fc;
	16'hb27 : data <= 32'h130e0011;
	16'hb28 : data <= 32'h13020000;
	16'hb29 : data <= 32'h97500000;
	16'hb2a : data <= 32'h93800036;
	16'hb2b : data <= 32'h83c11000;
	16'hb2c : data <= 32'h13000000;
	16'hb2d : data <= 32'h13000000;
	16'hb2e : data <= 32'h13830100;
	16'hb2f : data <= 32'h930e0000;
	16'hb30 : data <= 32'h6304d301;
	16'hb31 : data <= 32'h6f401059;
	16'hb32 : data <= 32'h13021200;
	16'hb33 : data <= 32'h93022000;
	16'hb34 : data <= 32'he31a52fc;
	16'hb35 : data <= 32'h130e1011;
	16'hb36 : data <= 32'h13020000;
	16'hb37 : data <= 32'h97500000;
	16'hb38 : data <= 32'h93809032;
	16'hb39 : data <= 32'h83c11000;
	16'hb3a : data <= 32'h930e000f;
	16'hb3b : data <= 32'h6384d101;
	16'hb3c : data <= 32'h6f405056;
	16'hb3d : data <= 32'h13021200;
	16'hb3e : data <= 32'h93022000;
	16'hb3f : data <= 32'he31052fe;
	16'hb40 : data <= 32'h130e2011;
	16'hb41 : data <= 32'h13020000;
	16'hb42 : data <= 32'h97500000;
	16'hb43 : data <= 32'h9380e02f;
	16'hb44 : data <= 32'h13000000;
	16'hb45 : data <= 32'h83c11000;
	16'hb46 : data <= 32'h930ef000;
	16'hb47 : data <= 32'h6384d101;
	16'hb48 : data <= 32'h6f405053;
	16'hb49 : data <= 32'h13021200;
	16'hb4a : data <= 32'h93022000;
	16'hb4b : data <= 32'he31e52fc;
	16'hb4c : data <= 32'h130e3011;
	16'hb4d : data <= 32'h13020000;
	16'hb4e : data <= 32'h97500000;
	16'hb4f : data <= 32'h9380c02c;
	16'hb50 : data <= 32'h13000000;
	16'hb51 : data <= 32'h13000000;
	16'hb52 : data <= 32'h83c11000;
	16'hb53 : data <= 32'h930e0000;
	16'hb54 : data <= 32'h6384d101;
	16'hb55 : data <= 32'h6f401050;
	16'hb56 : data <= 32'h13021200;
	16'hb57 : data <= 32'h93022000;
	16'hb58 : data <= 32'he31c52fc;
	16'hb59 : data <= 32'h97510000;
	16'hb5a : data <= 32'h9381012a;
	16'hb5b : data <= 32'h03c10100;
	16'hb5c : data <= 32'h13012000;
	16'hb5d : data <= 32'h930e2000;
	16'hb5e : data <= 32'h130e4011;
	16'hb5f : data <= 32'h6304d101;
	16'hb60 : data <= 32'h6f40504d;
	16'hb61 : data <= 32'h97510000;
	16'hb62 : data <= 32'h93810128;
	16'hb63 : data <= 32'h03c10100;
	16'hb64 : data <= 32'h13000000;
	16'hb65 : data <= 32'h13012000;
	16'hb66 : data <= 32'h930e2000;
	16'hb67 : data <= 32'h130e5011;
	16'hb68 : data <= 32'h6304d101;
	16'hb69 : data <= 32'h6f40104b;
	16'hb6a : data <= 32'h97500000;
	16'hb6b : data <= 32'h93800026;
	16'hb6c : data <= 32'h83910000;
	16'hb6d : data <= 32'h930ef00f;
	16'hb6e : data <= 32'h130e6011;
	16'hb6f : data <= 32'h6384d101;
	16'hb70 : data <= 32'h6f405049;
	16'hb71 : data <= 32'h97500000;
	16'hb72 : data <= 32'h93804024;
	16'hb73 : data <= 32'h83912000;
	16'hb74 : data <= 32'h930e00f0;
	16'hb75 : data <= 32'h130e7011;
	16'hb76 : data <= 32'h6384d101;
	16'hb77 : data <= 32'h6f409047;
	16'hb78 : data <= 32'h97500000;
	16'hb79 : data <= 32'h93808022;
	16'hb7a : data <= 32'h83914000;
	16'hb7b : data <= 32'hb71e0000;
	16'hb7c : data <= 32'h938e0eff;
	16'hb7d : data <= 32'h130e8011;
	16'hb7e : data <= 32'h6384d101;
	16'hb7f : data <= 32'h6f409045;
	16'hb80 : data <= 32'h97500000;
	16'hb81 : data <= 32'h93808020;
	16'hb82 : data <= 32'h83916000;
	16'hb83 : data <= 32'hb7feffff;
	16'hb84 : data <= 32'h938efe00;
	16'hb85 : data <= 32'h130e9011;
	16'hb86 : data <= 32'h6384d101;
	16'hb87 : data <= 32'h6f409043;
	16'hb88 : data <= 32'h97500000;
	16'hb89 : data <= 32'h9380e01e;
	16'hb8a : data <= 32'h8391a0ff;
	16'hb8b : data <= 32'h930ef00f;
	16'hb8c : data <= 32'h130ea011;
	16'hb8d : data <= 32'h6384d101;
	16'hb8e : data <= 32'h6f40d041;
	16'hb8f : data <= 32'h97500000;
	16'hb90 : data <= 32'h9380201d;
	16'hb91 : data <= 32'h8391c0ff;
	16'hb92 : data <= 32'h930e00f0;
	16'hb93 : data <= 32'h130eb011;
	16'hb94 : data <= 32'h6384d101;
	16'hb95 : data <= 32'h6f401040;
	16'hb96 : data <= 32'h97500000;
	16'hb97 : data <= 32'h9380601b;
	16'hb98 : data <= 32'h8391e0ff;
	16'hb99 : data <= 32'hb71e0000;
	16'hb9a : data <= 32'h938e0eff;
	16'hb9b : data <= 32'h130ec011;
	16'hb9c : data <= 32'h6384d101;
	16'hb9d : data <= 32'h6f40103e;
	16'hb9e : data <= 32'h97500000;
	16'hb9f : data <= 32'h93806019;
	16'hba0 : data <= 32'h83910000;
	16'hba1 : data <= 32'hb7feffff;
	16'hba2 : data <= 32'h938efe00;
	16'hba3 : data <= 32'h130ed011;
	16'hba4 : data <= 32'h6384d101;
	16'hba5 : data <= 32'h6f40103c;
	16'hba6 : data <= 32'h97500000;
	16'hba7 : data <= 32'h93800017;
	16'hba8 : data <= 32'h938000fe;
	16'hba9 : data <= 32'h83910002;
	16'hbaa : data <= 32'h930ef00f;
	16'hbab : data <= 32'h130ee011;
	16'hbac : data <= 32'h6384d101;
	16'hbad : data <= 32'h6f40103a;
	16'hbae : data <= 32'h97500000;
	16'hbaf : data <= 32'h93800015;
	16'hbb0 : data <= 32'h9380b0ff;
	16'hbb1 : data <= 32'h83917000;
	16'hbb2 : data <= 32'h930e00f0;
	16'hbb3 : data <= 32'h130ef011;
	16'hbb4 : data <= 32'h6384d101;
	16'hbb5 : data <= 32'h6f401038;
	16'hbb6 : data <= 32'h130e0012;
	16'hbb7 : data <= 32'h13020000;
	16'hbb8 : data <= 32'h97500000;
	16'hbb9 : data <= 32'h9380a012;
	16'hbba : data <= 32'h83912000;
	16'hbbb : data <= 32'h13830100;
	16'hbbc : data <= 32'hb71e0000;
	16'hbbd : data <= 32'h938e0eff;
	16'hbbe : data <= 32'h6304d301;
	16'hbbf : data <= 32'h6f409035;
	16'hbc0 : data <= 32'h13021200;
	16'hbc1 : data <= 32'h93022000;
	16'hbc2 : data <= 32'he31c52fc;
	16'hbc3 : data <= 32'h130e1012;
	16'hbc4 : data <= 32'h13020000;
	16'hbc5 : data <= 32'h97500000;
	16'hbc6 : data <= 32'h9380800f;
	16'hbc7 : data <= 32'h83912000;
	16'hbc8 : data <= 32'h13000000;
	16'hbc9 : data <= 32'h13830100;
	16'hbca : data <= 32'hb7feffff;
	16'hbcb : data <= 32'h938efe00;
	16'hbcc : data <= 32'h6304d301;
	16'hbcd : data <= 32'h6f401032;
	16'hbce : data <= 32'h13021200;
	16'hbcf : data <= 32'h93022000;
	16'hbd0 : data <= 32'he31a52fc;
	16'hbd1 : data <= 32'h130e2012;
	16'hbd2 : data <= 32'h13020000;
	16'hbd3 : data <= 32'h97500000;
	16'hbd4 : data <= 32'h9380c00b;
	16'hbd5 : data <= 32'h83912000;
	16'hbd6 : data <= 32'h13000000;
	16'hbd7 : data <= 32'h13000000;
	16'hbd8 : data <= 32'h13830100;
	16'hbd9 : data <= 32'h930e00f0;
	16'hbda : data <= 32'h6304d301;
	16'hbdb : data <= 32'h6f40902e;
	16'hbdc : data <= 32'h13021200;
	16'hbdd : data <= 32'h93022000;
	16'hbde : data <= 32'he31a52fc;
	16'hbdf : data <= 32'h130e3012;
	16'hbe0 : data <= 32'h13020000;
	16'hbe1 : data <= 32'h97500000;
	16'hbe2 : data <= 32'h93806008;
	16'hbe3 : data <= 32'h83912000;
	16'hbe4 : data <= 32'hb71e0000;
	16'hbe5 : data <= 32'h938e0eff;
	16'hbe6 : data <= 32'h6384d101;
	16'hbe7 : data <= 32'h6f40902b;
	16'hbe8 : data <= 32'h13021200;
	16'hbe9 : data <= 32'h93022000;
	16'hbea : data <= 32'he31e52fc;
	16'hbeb : data <= 32'h130e4012;
	16'hbec : data <= 32'h13020000;
	16'hbed : data <= 32'h97500000;
	16'hbee : data <= 32'h93808005;
	16'hbef : data <= 32'h13000000;
	16'hbf0 : data <= 32'h83912000;
	16'hbf1 : data <= 32'hb7feffff;
	16'hbf2 : data <= 32'h938efe00;
	16'hbf3 : data <= 32'h6384d101;
	16'hbf4 : data <= 32'h6f405028;
	16'hbf5 : data <= 32'h13021200;
	16'hbf6 : data <= 32'h93022000;
	16'hbf7 : data <= 32'he31c52fc;
	16'hbf8 : data <= 32'h130e5012;
	16'hbf9 : data <= 32'h13020000;
	16'hbfa : data <= 32'h97500000;
	16'hbfb : data <= 32'h93800002;
	16'hbfc : data <= 32'h13000000;
	16'hbfd : data <= 32'h13000000;
	16'hbfe : data <= 32'h83912000;
	16'hbff : data <= 32'h930e00f0;
	16'hc00 : data <= 32'h6384d101;
	16'hc01 : data <= 32'h6f401025;
	16'hc02 : data <= 32'h13021200;
	16'hc03 : data <= 32'h93022000;
	16'hc04 : data <= 32'he31c52fc;
	16'hc05 : data <= 32'h97510000;
	16'hc06 : data <= 32'h938141ff;
	16'hc07 : data <= 32'h03910100;
	16'hc08 : data <= 32'h13012000;
	16'hc09 : data <= 32'h930e2000;
	16'hc0a : data <= 32'h130e6012;
	16'hc0b : data <= 32'h6304d101;
	16'hc0c : data <= 32'h6f405022;
	16'hc0d : data <= 32'h97510000;
	16'hc0e : data <= 32'h938141fd;
	16'hc0f : data <= 32'h03910100;
	16'hc10 : data <= 32'h13000000;
	16'hc11 : data <= 32'h13012000;
	16'hc12 : data <= 32'h930e2000;
	16'hc13 : data <= 32'h130e7012;
	16'hc14 : data <= 32'h6304d101;
	16'hc15 : data <= 32'h6f401020;
	16'hc16 : data <= 32'h97500000;
	16'hc17 : data <= 32'h938080fb;
	16'hc18 : data <= 32'h83d10000;
	16'hc19 : data <= 32'h930ef00f;
	16'hc1a : data <= 32'h130e8012;
	16'hc1b : data <= 32'h6384d101;
	16'hc1c : data <= 32'h6f40501e;
	16'hc1d : data <= 32'h97500000;
	16'hc1e : data <= 32'h9380c0f9;
	16'hc1f : data <= 32'h83d12000;
	16'hc20 : data <= 32'hb70e0100;
	16'hc21 : data <= 32'h938e0ef0;
	16'hc22 : data <= 32'h130e9012;
	16'hc23 : data <= 32'h6384d101;
	16'hc24 : data <= 32'h6f40501c;
	16'hc25 : data <= 32'h97500000;
	16'hc26 : data <= 32'h9380c0f7;
	16'hc27 : data <= 32'h83d14000;
	16'hc28 : data <= 32'hb71e0000;
	16'hc29 : data <= 32'h938e0eff;
	16'hc2a : data <= 32'h130ea012;
	16'hc2b : data <= 32'h6384d101;
	16'hc2c : data <= 32'h6f40501a;
	16'hc2d : data <= 32'h97500000;
	16'hc2e : data <= 32'h9380c0f5;
	16'hc2f : data <= 32'h83d16000;
	16'hc30 : data <= 32'hb7fe0000;
	16'hc31 : data <= 32'h938efe00;
	16'hc32 : data <= 32'h130eb012;
	16'hc33 : data <= 32'h6384d101;
	16'hc34 : data <= 32'h6f405018;
	16'hc35 : data <= 32'h97500000;
	16'hc36 : data <= 32'h938020f4;
	16'hc37 : data <= 32'h83d1a0ff;
	16'hc38 : data <= 32'h930ef00f;
	16'hc39 : data <= 32'h130ec012;
	16'hc3a : data <= 32'h6384d101;
	16'hc3b : data <= 32'h6f409016;
	16'hc3c : data <= 32'h97500000;
	16'hc3d : data <= 32'h938060f2;
	16'hc3e : data <= 32'h83d1c0ff;
	16'hc3f : data <= 32'hb70e0100;
	16'hc40 : data <= 32'h938e0ef0;
	16'hc41 : data <= 32'h130ed012;
	16'hc42 : data <= 32'h6384d101;
	16'hc43 : data <= 32'h6f409014;
	16'hc44 : data <= 32'h97500000;
	16'hc45 : data <= 32'h938060f0;
	16'hc46 : data <= 32'h83d1e0ff;
	16'hc47 : data <= 32'hb71e0000;
	16'hc48 : data <= 32'h938e0eff;
	16'hc49 : data <= 32'h130ee012;
	16'hc4a : data <= 32'h6384d101;
	16'hc4b : data <= 32'h6f409012;
	16'hc4c : data <= 32'h97500000;
	16'hc4d : data <= 32'h938060ee;
	16'hc4e : data <= 32'h83d10000;
	16'hc4f : data <= 32'hb7fe0000;
	16'hc50 : data <= 32'h938efe00;
	16'hc51 : data <= 32'h130ef012;
	16'hc52 : data <= 32'h6384d101;
	16'hc53 : data <= 32'h6f409010;
	16'hc54 : data <= 32'h97500000;
	16'hc55 : data <= 32'h938000ec;
	16'hc56 : data <= 32'h938000fe;
	16'hc57 : data <= 32'h83d10002;
	16'hc58 : data <= 32'h930ef00f;
	16'hc59 : data <= 32'h130e0013;
	16'hc5a : data <= 32'h6384d101;
	16'hc5b : data <= 32'h6f40900e;
	16'hc5c : data <= 32'h97500000;
	16'hc5d : data <= 32'h938000ea;
	16'hc5e : data <= 32'h9380b0ff;
	16'hc5f : data <= 32'h83d17000;
	16'hc60 : data <= 32'hb70e0100;
	16'hc61 : data <= 32'h938e0ef0;
	16'hc62 : data <= 32'h130e1013;
	16'hc63 : data <= 32'h6384d101;
	16'hc64 : data <= 32'h6f40500c;
	16'hc65 : data <= 32'h130e2013;
	16'hc66 : data <= 32'h13020000;
	16'hc67 : data <= 32'h97500000;
	16'hc68 : data <= 32'h938060e7;
	16'hc69 : data <= 32'h83d12000;
	16'hc6a : data <= 32'h13830100;
	16'hc6b : data <= 32'hb71e0000;
	16'hc6c : data <= 32'h938e0eff;
	16'hc6d : data <= 32'h6304d301;
	16'hc6e : data <= 32'h6f40d009;
	16'hc6f : data <= 32'h13021200;
	16'hc70 : data <= 32'h93022000;
	16'hc71 : data <= 32'he31c52fc;
	16'hc72 : data <= 32'h130e3013;
	16'hc73 : data <= 32'h13020000;
	16'hc74 : data <= 32'h97500000;
	16'hc75 : data <= 32'h938040e4;
	16'hc76 : data <= 32'h83d12000;
	16'hc77 : data <= 32'h13000000;
	16'hc78 : data <= 32'h13830100;
	16'hc79 : data <= 32'hb7fe0000;
	16'hc7a : data <= 32'h938efe00;
	16'hc7b : data <= 32'h6304d301;
	16'hc7c : data <= 32'h6f405006;
	16'hc7d : data <= 32'h13021200;
	16'hc7e : data <= 32'h93022000;
	16'hc7f : data <= 32'he31a52fc;
	16'hc80 : data <= 32'h130e4013;
	16'hc81 : data <= 32'h13020000;
	16'hc82 : data <= 32'h97500000;
	16'hc83 : data <= 32'h938080e0;
	16'hc84 : data <= 32'h83d12000;
	16'hc85 : data <= 32'h13000000;
	16'hc86 : data <= 32'h13000000;
	16'hc87 : data <= 32'h13830100;
	16'hc88 : data <= 32'hb70e0100;
	16'hc89 : data <= 32'h938e0ef0;
	16'hc8a : data <= 32'h6304d301;
	16'hc8b : data <= 32'h6f409002;
	16'hc8c : data <= 32'h13021200;
	16'hc8d : data <= 32'h93022000;
	16'hc8e : data <= 32'he31852fc;
	16'hc8f : data <= 32'h130e5013;
	16'hc90 : data <= 32'h13020000;
	16'hc91 : data <= 32'h97500000;
	16'hc92 : data <= 32'h9380e0dc;
	16'hc93 : data <= 32'h83d12000;
	16'hc94 : data <= 32'hb71e0000;
	16'hc95 : data <= 32'h938e0eff;
	16'hc96 : data <= 32'h6384d101;
	16'hc97 : data <= 32'h6f40807f;
	16'hc98 : data <= 32'h13021200;
	16'hc99 : data <= 32'h93022000;
	16'hc9a : data <= 32'he31e52fc;
	16'hc9b : data <= 32'h130e6013;
	16'hc9c : data <= 32'h13020000;
	16'hc9d : data <= 32'h97500000;
	16'hc9e : data <= 32'h938000da;
	16'hc9f : data <= 32'h13000000;
	16'hca0 : data <= 32'h83d12000;
	16'hca1 : data <= 32'hb7fe0000;
	16'hca2 : data <= 32'h938efe00;
	16'hca3 : data <= 32'h6384d101;
	16'hca4 : data <= 32'h6f40407c;
	16'hca5 : data <= 32'h13021200;
	16'hca6 : data <= 32'h93022000;
	16'hca7 : data <= 32'he31c52fc;
	16'hca8 : data <= 32'h130e7013;
	16'hca9 : data <= 32'h13020000;
	16'hcaa : data <= 32'h97500000;
	16'hcab : data <= 32'h938080d6;
	16'hcac : data <= 32'h13000000;
	16'hcad : data <= 32'h13000000;
	16'hcae : data <= 32'h83d12000;
	16'hcaf : data <= 32'hb70e0100;
	16'hcb0 : data <= 32'h938e0ef0;
	16'hcb1 : data <= 32'h6384d101;
	16'hcb2 : data <= 32'h6f40c078;
	16'hcb3 : data <= 32'h13021200;
	16'hcb4 : data <= 32'h93022000;
	16'hcb5 : data <= 32'he31a52fc;
	16'hcb6 : data <= 32'h97510000;
	16'hcb7 : data <= 32'h938181d3;
	16'hcb8 : data <= 32'h03d10100;
	16'hcb9 : data <= 32'h13012000;
	16'hcba : data <= 32'h930e2000;
	16'hcbb : data <= 32'h130e8013;
	16'hcbc : data <= 32'h6304d101;
	16'hcbd : data <= 32'h6f400076;
	16'hcbe : data <= 32'h97510000;
	16'hcbf : data <= 32'h938181d1;
	16'hcc0 : data <= 32'h03d10100;
	16'hcc1 : data <= 32'h13000000;
	16'hcc2 : data <= 32'h13012000;
	16'hcc3 : data <= 32'h930e2000;
	16'hcc4 : data <= 32'h130e9013;
	16'hcc5 : data <= 32'h6304d101;
	16'hcc6 : data <= 32'h6f40c073;
	16'hcc7 : data <= 32'hb7000000;
	16'hcc8 : data <= 32'h930e0000;
	16'hcc9 : data <= 32'h130ea013;
	16'hcca : data <= 32'h6384d001;
	16'hccb : data <= 32'h6f408072;
	16'hccc : data <= 32'hb7f0ffff;
	16'hccd : data <= 32'h93d01040;
	16'hcce : data <= 32'h930e0080;
	16'hccf : data <= 32'h130eb013;
	16'hcd0 : data <= 32'h6384d001;
	16'hcd1 : data <= 32'h6f400071;
	16'hcd2 : data <= 32'hb7f0ff7f;
	16'hcd3 : data <= 32'h93d04041;
	16'hcd4 : data <= 32'h930ef07f;
	16'hcd5 : data <= 32'h130ec013;
	16'hcd6 : data <= 32'h6384d001;
	16'hcd7 : data <= 32'h6f40806f;
	16'hcd8 : data <= 32'hb7000080;
	16'hcd9 : data <= 32'h93d04041;
	16'hcda : data <= 32'h930e0080;
	16'hcdb : data <= 32'h130ed013;
	16'hcdc : data <= 32'h6384d001;
	16'hcdd : data <= 32'h6f40006e;
	16'hcde : data <= 32'h37000080;
	16'hcdf : data <= 32'h930e0000;
	16'hce0 : data <= 32'h130ee013;
	16'hce1 : data <= 32'h6304d001;
	16'hce2 : data <= 32'h6f40c06c;
	16'hce3 : data <= 32'h97500000;
	16'hce4 : data <= 32'h9380c0c8;
	16'hce5 : data <= 32'h83a10000;
	16'hce6 : data <= 32'hb70eff00;
	16'hce7 : data <= 32'h938efe0f;
	16'hce8 : data <= 32'h130ef013;
	16'hce9 : data <= 32'h6384d101;
	16'hcea : data <= 32'h6f40c06a;
	16'hceb : data <= 32'h97500000;
	16'hcec : data <= 32'h9380c0c6;
	16'hced : data <= 32'h83a14000;
	16'hcee : data <= 32'hb70e01ff;
	16'hcef : data <= 32'h938e0ef0;
	16'hcf0 : data <= 32'h130e0014;
	16'hcf1 : data <= 32'h6384d101;
	16'hcf2 : data <= 32'h6f40c068;
	16'hcf3 : data <= 32'h97500000;
	16'hcf4 : data <= 32'h9380c0c4;
	16'hcf5 : data <= 32'h83a18000;
	16'hcf6 : data <= 32'hb71ef00f;
	16'hcf7 : data <= 32'h938e0eff;
	16'hcf8 : data <= 32'h130e1014;
	16'hcf9 : data <= 32'h6384d101;
	16'hcfa : data <= 32'h6f40c066;
	16'hcfb : data <= 32'h97500000;
	16'hcfc : data <= 32'h9380c0c2;
	16'hcfd : data <= 32'h83a1c000;
	16'hcfe : data <= 32'hb7fe0ff0;
	16'hcff : data <= 32'h938efe00;
	16'hd00 : data <= 32'h130e2014;
	16'hd01 : data <= 32'h6384d101;
	16'hd02 : data <= 32'h6f40c064;
	16'hd03 : data <= 32'h97500000;
	16'hd04 : data <= 32'h938080c1;
	16'hd05 : data <= 32'h83a140ff;
	16'hd06 : data <= 32'hb70eff00;
	16'hd07 : data <= 32'h938efe0f;
	16'hd08 : data <= 32'h130e3014;
	16'hd09 : data <= 32'h6384d101;
	16'hd0a : data <= 32'h6f40c062;
	16'hd0b : data <= 32'h97500000;
	16'hd0c : data <= 32'h938080bf;
	16'hd0d : data <= 32'h83a180ff;
	16'hd0e : data <= 32'hb70e01ff;
	16'hd0f : data <= 32'h938e0ef0;
	16'hd10 : data <= 32'h130e4014;
	16'hd11 : data <= 32'h6384d101;
	16'hd12 : data <= 32'h6f40c060;
	16'hd13 : data <= 32'h97500000;
	16'hd14 : data <= 32'h938080bd;
	16'hd15 : data <= 32'h83a1c0ff;
	16'hd16 : data <= 32'hb71ef00f;
	16'hd17 : data <= 32'h938e0eff;
	16'hd18 : data <= 32'h130e5014;
	16'hd19 : data <= 32'h6384d101;
	16'hd1a : data <= 32'h6f40c05e;
	16'hd1b : data <= 32'h97500000;
	16'hd1c : data <= 32'h938080bb;
	16'hd1d : data <= 32'h83a10000;
	16'hd1e : data <= 32'hb7fe0ff0;
	16'hd1f : data <= 32'h938efe00;
	16'hd20 : data <= 32'h130e6014;
	16'hd21 : data <= 32'h6384d101;
	16'hd22 : data <= 32'h6f40c05c;
	16'hd23 : data <= 32'h97500000;
	16'hd24 : data <= 32'h9380c0b8;
	16'hd25 : data <= 32'h938000fe;
	16'hd26 : data <= 32'h83a10002;
	16'hd27 : data <= 32'hb70eff00;
	16'hd28 : data <= 32'h938efe0f;
	16'hd29 : data <= 32'h130e7014;
	16'hd2a : data <= 32'h6384d101;
	16'hd2b : data <= 32'h6f40805a;
	16'hd2c : data <= 32'h97500000;
	16'hd2d : data <= 32'h938080b6;
	16'hd2e : data <= 32'h9380d0ff;
	16'hd2f : data <= 32'h83a17000;
	16'hd30 : data <= 32'hb70e01ff;
	16'hd31 : data <= 32'h938e0ef0;
	16'hd32 : data <= 32'h130e8014;
	16'hd33 : data <= 32'h6384d101;
	16'hd34 : data <= 32'h6f404058;
	16'hd35 : data <= 32'h130e9014;
	16'hd36 : data <= 32'h13020000;
	16'hd37 : data <= 32'h97500000;
	16'hd38 : data <= 32'h938000b4;
	16'hd39 : data <= 32'h83a14000;
	16'hd3a : data <= 32'h13830100;
	16'hd3b : data <= 32'hb71ef00f;
	16'hd3c : data <= 32'h938e0eff;
	16'hd3d : data <= 32'h6304d301;
	16'hd3e : data <= 32'h6f40c055;
	16'hd3f : data <= 32'h13021200;
	16'hd40 : data <= 32'h93022000;
	16'hd41 : data <= 32'he31c52fc;
	16'hd42 : data <= 32'h130ea014;
	16'hd43 : data <= 32'h13020000;
	16'hd44 : data <= 32'h97500000;
	16'hd45 : data <= 32'h938000b1;
	16'hd46 : data <= 32'h83a14000;
	16'hd47 : data <= 32'h13000000;
	16'hd48 : data <= 32'h13830100;
	16'hd49 : data <= 32'hb7fe0ff0;
	16'hd4a : data <= 32'h938efe00;
	16'hd4b : data <= 32'h6304d301;
	16'hd4c : data <= 32'h6f404052;
	16'hd4d : data <= 32'h13021200;
	16'hd4e : data <= 32'h93022000;
	16'hd4f : data <= 32'he31a52fc;
	16'hd50 : data <= 32'h130eb014;
	16'hd51 : data <= 32'h13020000;
	16'hd52 : data <= 32'h97500000;
	16'hd53 : data <= 32'h938000ad;
	16'hd54 : data <= 32'h83a14000;
	16'hd55 : data <= 32'h13000000;
	16'hd56 : data <= 32'h13000000;
	16'hd57 : data <= 32'h13830100;
	16'hd58 : data <= 32'hb70e01ff;
	16'hd59 : data <= 32'h938e0ef0;
	16'hd5a : data <= 32'h6304d301;
	16'hd5b : data <= 32'h6f40804e;
	16'hd5c : data <= 32'h13021200;
	16'hd5d : data <= 32'h93022000;
	16'hd5e : data <= 32'he31852fc;
	16'hd5f : data <= 32'h130ec014;
	16'hd60 : data <= 32'h13020000;
	16'hd61 : data <= 32'h97500000;
	16'hd62 : data <= 32'h938080a9;
	16'hd63 : data <= 32'h83a14000;
	16'hd64 : data <= 32'hb71ef00f;
	16'hd65 : data <= 32'h938e0eff;
	16'hd66 : data <= 32'h6384d101;
	16'hd67 : data <= 32'h6f40804b;
	16'hd68 : data <= 32'h13021200;
	16'hd69 : data <= 32'h93022000;
	16'hd6a : data <= 32'he31e52fc;
	16'hd6b : data <= 32'h130ed014;
	16'hd6c : data <= 32'h13020000;
	16'hd6d : data <= 32'h97500000;
	16'hd6e : data <= 32'h9380c0a6;
	16'hd6f : data <= 32'h13000000;
	16'hd70 : data <= 32'h83a14000;
	16'hd71 : data <= 32'hb7fe0ff0;
	16'hd72 : data <= 32'h938efe00;
	16'hd73 : data <= 32'h6384d101;
	16'hd74 : data <= 32'h6f404048;
	16'hd75 : data <= 32'h13021200;
	16'hd76 : data <= 32'h93022000;
	16'hd77 : data <= 32'he31c52fc;
	16'hd78 : data <= 32'h130ee014;
	16'hd79 : data <= 32'h13020000;
	16'hd7a : data <= 32'h97500000;
	16'hd7b : data <= 32'h938000a3;
	16'hd7c : data <= 32'h13000000;
	16'hd7d : data <= 32'h13000000;
	16'hd7e : data <= 32'h83a14000;
	16'hd7f : data <= 32'hb70e01ff;
	16'hd80 : data <= 32'h938e0ef0;
	16'hd81 : data <= 32'h6384d101;
	16'hd82 : data <= 32'h6f40c044;
	16'hd83 : data <= 32'h13021200;
	16'hd84 : data <= 32'h93022000;
	16'hd85 : data <= 32'he31a52fc;
	16'hd86 : data <= 32'h97510000;
	16'hd87 : data <= 32'h938101a0;
	16'hd88 : data <= 32'h03a10100;
	16'hd89 : data <= 32'h13012000;
	16'hd8a : data <= 32'h930e2000;
	16'hd8b : data <= 32'h130ef014;
	16'hd8c : data <= 32'h6304d101;
	16'hd8d : data <= 32'h6f400042;
	16'hd8e : data <= 32'h97510000;
	16'hd8f : data <= 32'h9381019e;
	16'hd90 : data <= 32'h03a10100;
	16'hd91 : data <= 32'h13000000;
	16'hd92 : data <= 32'h13012000;
	16'hd93 : data <= 32'h930e2000;
	16'hd94 : data <= 32'h130e0015;
	16'hd95 : data <= 32'h6304d101;
	16'hd96 : data <= 32'h6f40c03f;
	16'hd97 : data <= 32'hb70001ff;
	16'hd98 : data <= 32'h938000f0;
	16'hd99 : data <= 32'h37110f0f;
	16'hd9a : data <= 32'h1301f1f0;
	16'hd9b : data <= 32'hb3e12000;
	16'hd9c : data <= 32'hb70e10ff;
	16'hd9d : data <= 32'h938efef0;
	16'hd9e : data <= 32'h130e1015;
	16'hd9f : data <= 32'h6384d101;
	16'hda0 : data <= 32'h6f40403d;
	16'hda1 : data <= 32'hb710f00f;
	16'hda2 : data <= 32'h938000ff;
	16'hda3 : data <= 32'h37f1f0f0;
	16'hda4 : data <= 32'h1301010f;
	16'hda5 : data <= 32'hb3e12000;
	16'hda6 : data <= 32'hb70ef1ff;
	16'hda7 : data <= 32'h938e0eff;
	16'hda8 : data <= 32'h130e2015;
	16'hda9 : data <= 32'h6384d101;
	16'hdaa : data <= 32'h6f40c03a;
	16'hdab : data <= 32'hb700ff00;
	16'hdac : data <= 32'h9380f00f;
	16'hdad : data <= 32'h37110f0f;
	16'hdae : data <= 32'h1301f1f0;
	16'hdaf : data <= 32'hb3e12000;
	16'hdb0 : data <= 32'hb71eff0f;
	16'hdb1 : data <= 32'h938efeff;
	16'hdb2 : data <= 32'h130e3015;
	16'hdb3 : data <= 32'h6384d101;
	16'hdb4 : data <= 32'h6f404038;
	16'hdb5 : data <= 32'hb7f00ff0;
	16'hdb6 : data <= 32'h9380f000;
	16'hdb7 : data <= 32'h37f1f0f0;
	16'hdb8 : data <= 32'h1301010f;
	16'hdb9 : data <= 32'hb3e12000;
	16'hdba : data <= 32'hb7fefff0;
	16'hdbb : data <= 32'h938efe0f;
	16'hdbc : data <= 32'h130e4015;
	16'hdbd : data <= 32'h6384d101;
	16'hdbe : data <= 32'h6f40c035;
	16'hdbf : data <= 32'hb70001ff;
	16'hdc0 : data <= 32'h938000f0;
	16'hdc1 : data <= 32'h37110f0f;
	16'hdc2 : data <= 32'h1301f1f0;
	16'hdc3 : data <= 32'hb3e02000;
	16'hdc4 : data <= 32'hb70e10ff;
	16'hdc5 : data <= 32'h938efef0;
	16'hdc6 : data <= 32'h130e5015;
	16'hdc7 : data <= 32'h6384d001;
	16'hdc8 : data <= 32'h6f404033;
	16'hdc9 : data <= 32'hb70001ff;
	16'hdca : data <= 32'h938000f0;
	16'hdcb : data <= 32'h37110f0f;
	16'hdcc : data <= 32'h1301f1f0;
	16'hdcd : data <= 32'h33e12000;
	16'hdce : data <= 32'hb70e10ff;
	16'hdcf : data <= 32'h938efef0;
	16'hdd0 : data <= 32'h130e6015;
	16'hdd1 : data <= 32'h6304d101;
	16'hdd2 : data <= 32'h6f40c030;
	16'hdd3 : data <= 32'hb70001ff;
	16'hdd4 : data <= 32'h938000f0;
	16'hdd5 : data <= 32'hb3e01000;
	16'hdd6 : data <= 32'hb70e01ff;
	16'hdd7 : data <= 32'h938e0ef0;
	16'hdd8 : data <= 32'h130e7015;
	16'hdd9 : data <= 32'h6384d001;
	16'hdda : data <= 32'h6f40c02e;
	16'hddb : data <= 32'h13020000;
	16'hddc : data <= 32'hb70001ff;
	16'hddd : data <= 32'h938000f0;
	16'hdde : data <= 32'h37110f0f;
	16'hddf : data <= 32'h1301f1f0;
	16'hde0 : data <= 32'hb3e12000;
	16'hde1 : data <= 32'h13830100;
	16'hde2 : data <= 32'h13021200;
	16'hde3 : data <= 32'h93022000;
	16'hde4 : data <= 32'he31052fe;
	16'hde5 : data <= 32'hb70e10ff;
	16'hde6 : data <= 32'h938efef0;
	16'hde7 : data <= 32'h130e8015;
	16'hde8 : data <= 32'h6304d301;
	16'hde9 : data <= 32'h6f40002b;
	16'hdea : data <= 32'h13020000;
	16'hdeb : data <= 32'hb710f00f;
	16'hdec : data <= 32'h938000ff;
	16'hded : data <= 32'h37f1f0f0;
	16'hdee : data <= 32'h1301010f;
	16'hdef : data <= 32'hb3e12000;
	16'hdf0 : data <= 32'h13000000;
	16'hdf1 : data <= 32'h13830100;
	16'hdf2 : data <= 32'h13021200;
	16'hdf3 : data <= 32'h93022000;
	16'hdf4 : data <= 32'he31e52fc;
	16'hdf5 : data <= 32'hb70ef1ff;
	16'hdf6 : data <= 32'h938e0eff;
	16'hdf7 : data <= 32'h130e9015;
	16'hdf8 : data <= 32'h6304d301;
	16'hdf9 : data <= 32'h6f400027;
	16'hdfa : data <= 32'h13020000;
	16'hdfb : data <= 32'hb700ff00;
	16'hdfc : data <= 32'h9380f00f;
	16'hdfd : data <= 32'h37110f0f;
	16'hdfe : data <= 32'h1301f1f0;
	16'hdff : data <= 32'hb3e12000;
	16'he00 : data <= 32'h13000000;
	16'he01 : data <= 32'h13000000;
	16'he02 : data <= 32'h13830100;
	16'he03 : data <= 32'h13021200;
	16'he04 : data <= 32'h93022000;
	16'he05 : data <= 32'he31c52fc;
	16'he06 : data <= 32'hb71eff0f;
	16'he07 : data <= 32'h938efeff;
	16'he08 : data <= 32'h130ea015;
	16'he09 : data <= 32'h6304d301;
	16'he0a : data <= 32'h6f40c022;
	16'he0b : data <= 32'h13020000;
	16'he0c : data <= 32'hb70001ff;
	16'he0d : data <= 32'h938000f0;
	16'he0e : data <= 32'h37110f0f;
	16'he0f : data <= 32'h1301f1f0;
	16'he10 : data <= 32'hb3e12000;
	16'he11 : data <= 32'h13021200;
	16'he12 : data <= 32'h93022000;
	16'he13 : data <= 32'he31252fe;
	16'he14 : data <= 32'hb70e10ff;
	16'he15 : data <= 32'h938efef0;
	16'he16 : data <= 32'h130eb015;
	16'he17 : data <= 32'h6384d101;
	16'he18 : data <= 32'h6f40401f;
	16'he19 : data <= 32'h13020000;
	16'he1a : data <= 32'hb710f00f;
	16'he1b : data <= 32'h938000ff;
	16'he1c : data <= 32'h37f1f0f0;
	16'he1d : data <= 32'h1301010f;
	16'he1e : data <= 32'h13000000;
	16'he1f : data <= 32'hb3e12000;
	16'he20 : data <= 32'h13021200;
	16'he21 : data <= 32'h93022000;
	16'he22 : data <= 32'he31052fe;
	16'he23 : data <= 32'hb70ef1ff;
	16'he24 : data <= 32'h938e0eff;
	16'he25 : data <= 32'h130ec015;
	16'he26 : data <= 32'h6384d101;
	16'he27 : data <= 32'h6f40801b;
	16'he28 : data <= 32'h13020000;
	16'he29 : data <= 32'hb700ff00;
	16'he2a : data <= 32'h9380f00f;
	16'he2b : data <= 32'h37110f0f;
	16'he2c : data <= 32'h1301f1f0;
	16'he2d : data <= 32'h13000000;
	16'he2e : data <= 32'h13000000;
	16'he2f : data <= 32'hb3e12000;
	16'he30 : data <= 32'h13021200;
	16'he31 : data <= 32'h93022000;
	16'he32 : data <= 32'he31e52fc;
	16'he33 : data <= 32'hb71eff0f;
	16'he34 : data <= 32'h938efeff;
	16'he35 : data <= 32'h130ed015;
	16'he36 : data <= 32'h6384d101;
	16'he37 : data <= 32'h6f408017;
	16'he38 : data <= 32'h13020000;
	16'he39 : data <= 32'hb70001ff;
	16'he3a : data <= 32'h938000f0;
	16'he3b : data <= 32'h13000000;
	16'he3c : data <= 32'h37110f0f;
	16'he3d : data <= 32'h1301f1f0;
	16'he3e : data <= 32'hb3e12000;
	16'he3f : data <= 32'h13021200;
	16'he40 : data <= 32'h93022000;
	16'he41 : data <= 32'he31052fe;
	16'he42 : data <= 32'hb70e10ff;
	16'he43 : data <= 32'h938efef0;
	16'he44 : data <= 32'h130ee015;
	16'he45 : data <= 32'h6384d101;
	16'he46 : data <= 32'h6f40c013;
	16'he47 : data <= 32'h13020000;
	16'he48 : data <= 32'hb710f00f;
	16'he49 : data <= 32'h938000ff;
	16'he4a : data <= 32'h13000000;
	16'he4b : data <= 32'h37f1f0f0;
	16'he4c : data <= 32'h1301010f;
	16'he4d : data <= 32'h13000000;
	16'he4e : data <= 32'hb3e12000;
	16'he4f : data <= 32'h13021200;
	16'he50 : data <= 32'h93022000;
	16'he51 : data <= 32'he31e52fc;
	16'he52 : data <= 32'hb70ef1ff;
	16'he53 : data <= 32'h938e0eff;
	16'he54 : data <= 32'h130ef015;
	16'he55 : data <= 32'h6384d101;
	16'he56 : data <= 32'h6f40c00f;
	16'he57 : data <= 32'h13020000;
	16'he58 : data <= 32'hb700ff00;
	16'he59 : data <= 32'h9380f00f;
	16'he5a : data <= 32'h13000000;
	16'he5b : data <= 32'h13000000;
	16'he5c : data <= 32'h37110f0f;
	16'he5d : data <= 32'h1301f1f0;
	16'he5e : data <= 32'hb3e12000;
	16'he5f : data <= 32'h13021200;
	16'he60 : data <= 32'h93022000;
	16'he61 : data <= 32'he31e52fc;
	16'he62 : data <= 32'hb71eff0f;
	16'he63 : data <= 32'h938efeff;
	16'he64 : data <= 32'h130e0016;
	16'he65 : data <= 32'h6384d101;
	16'he66 : data <= 32'h6f40c00b;
	16'he67 : data <= 32'h13020000;
	16'he68 : data <= 32'h37110f0f;
	16'he69 : data <= 32'h1301f1f0;
	16'he6a : data <= 32'hb70001ff;
	16'he6b : data <= 32'h938000f0;
	16'he6c : data <= 32'hb3e12000;
	16'he6d : data <= 32'h13021200;
	16'he6e : data <= 32'h93022000;
	16'he6f : data <= 32'he31252fe;
	16'he70 : data <= 32'hb70e10ff;
	16'he71 : data <= 32'h938efef0;
	16'he72 : data <= 32'h130e1016;
	16'he73 : data <= 32'h6384d101;
	16'he74 : data <= 32'h6f404008;
	16'he75 : data <= 32'h13020000;
	16'he76 : data <= 32'h37f1f0f0;
	16'he77 : data <= 32'h1301010f;
	16'he78 : data <= 32'hb710f00f;
	16'he79 : data <= 32'h938000ff;
	16'he7a : data <= 32'h13000000;
	16'he7b : data <= 32'hb3e12000;
	16'he7c : data <= 32'h13021200;
	16'he7d : data <= 32'h93022000;
	16'he7e : data <= 32'he31052fe;
	16'he7f : data <= 32'hb70ef1ff;
	16'he80 : data <= 32'h938e0eff;
	16'he81 : data <= 32'h130e2016;
	16'he82 : data <= 32'h6384d101;
	16'he83 : data <= 32'h6f408004;
	16'he84 : data <= 32'h13020000;
	16'he85 : data <= 32'h37110f0f;
	16'he86 : data <= 32'h1301f1f0;
	16'he87 : data <= 32'hb700ff00;
	16'he88 : data <= 32'h9380f00f;
	16'he89 : data <= 32'h13000000;
	16'he8a : data <= 32'h13000000;
	16'he8b : data <= 32'hb3e12000;
	16'he8c : data <= 32'h13021200;
	16'he8d : data <= 32'h93022000;
	16'he8e : data <= 32'he31e52fc;
	16'he8f : data <= 32'hb71eff0f;
	16'he90 : data <= 32'h938efeff;
	16'he91 : data <= 32'h130e3016;
	16'he92 : data <= 32'h6384d101;
	16'he93 : data <= 32'h6f408000;
	16'he94 : data <= 32'h13020000;
	16'he95 : data <= 32'h37110f0f;
	16'he96 : data <= 32'h1301f1f0;
	16'he97 : data <= 32'h13000000;
	16'he98 : data <= 32'hb70001ff;
	16'he99 : data <= 32'h938000f0;
	16'he9a : data <= 32'hb3e12000;
	16'he9b : data <= 32'h13021200;
	16'he9c : data <= 32'h93022000;
	16'he9d : data <= 32'he31052fe;
	16'he9e : data <= 32'hb70e10ff;
	16'he9f : data <= 32'h938efef0;
	16'hea0 : data <= 32'h130e4016;
	16'hea1 : data <= 32'h6384d101;
	16'hea2 : data <= 32'h6f30d07c;
	16'hea3 : data <= 32'h13020000;
	16'hea4 : data <= 32'h37f1f0f0;
	16'hea5 : data <= 32'h1301010f;
	16'hea6 : data <= 32'h13000000;
	16'hea7 : data <= 32'hb710f00f;
	16'hea8 : data <= 32'h938000ff;
	16'hea9 : data <= 32'h13000000;
	16'heaa : data <= 32'hb3e12000;
	16'heab : data <= 32'h13021200;
	16'heac : data <= 32'h93022000;
	16'head : data <= 32'he31e52fc;
	16'heae : data <= 32'hb70ef1ff;
	16'heaf : data <= 32'h938e0eff;
	16'heb0 : data <= 32'h130e5016;
	16'heb1 : data <= 32'h6384d101;
	16'heb2 : data <= 32'h6f30d078;
	16'heb3 : data <= 32'h13020000;
	16'heb4 : data <= 32'h37110f0f;
	16'heb5 : data <= 32'h1301f1f0;
	16'heb6 : data <= 32'h13000000;
	16'heb7 : data <= 32'h13000000;
	16'heb8 : data <= 32'hb700ff00;
	16'heb9 : data <= 32'h9380f00f;
	16'heba : data <= 32'hb3e12000;
	16'hebb : data <= 32'h13021200;
	16'hebc : data <= 32'h93022000;
	16'hebd : data <= 32'he31e52fc;
	16'hebe : data <= 32'hb71eff0f;
	16'hebf : data <= 32'h938efeff;
	16'hec0 : data <= 32'h130e6016;
	16'hec1 : data <= 32'h6384d101;
	16'hec2 : data <= 32'h6f30d074;
	16'hec3 : data <= 32'hb70001ff;
	16'hec4 : data <= 32'h938000f0;
	16'hec5 : data <= 32'h33611000;
	16'hec6 : data <= 32'hb70e01ff;
	16'hec7 : data <= 32'h938e0ef0;
	16'hec8 : data <= 32'h130e7016;
	16'hec9 : data <= 32'h6304d101;
	16'heca : data <= 32'h6f30d072;
	16'hecb : data <= 32'hb700ff00;
	16'hecc : data <= 32'h9380f00f;
	16'hecd : data <= 32'h33e10000;
	16'hece : data <= 32'hb70eff00;
	16'hecf : data <= 32'h938efe0f;
	16'hed0 : data <= 32'h130e8016;
	16'hed1 : data <= 32'h6304d101;
	16'hed2 : data <= 32'h6f30d070;
	16'hed3 : data <= 32'hb3600000;
	16'hed4 : data <= 32'h930e0000;
	16'hed5 : data <= 32'h130e9016;
	16'hed6 : data <= 32'h6384d001;
	16'hed7 : data <= 32'h6f30906f;
	16'hed8 : data <= 32'hb7101111;
	16'hed9 : data <= 32'h93801011;
	16'heda : data <= 32'h37212222;
	16'hedb : data <= 32'h13012122;
	16'hedc : data <= 32'h33e02000;
	16'hedd : data <= 32'h930e0000;
	16'hede : data <= 32'h130ea016;
	16'hedf : data <= 32'h6304d001;
	16'hee0 : data <= 32'h6f30506d;
	16'hee1 : data <= 32'hb70001ff;
	16'hee2 : data <= 32'h938000f0;
	16'hee3 : data <= 32'h93e1f0f0;
	16'hee4 : data <= 32'h930ef0f0;
	16'hee5 : data <= 32'h130eb016;
	16'hee6 : data <= 32'h6384d101;
	16'hee7 : data <= 32'h6f30906b;
	16'hee8 : data <= 32'hb710f00f;
	16'hee9 : data <= 32'h938000ff;
	16'heea : data <= 32'h93e1000f;
	16'heeb : data <= 32'hb71ef00f;
	16'heec : data <= 32'h938e0eff;
	16'heed : data <= 32'h130ec016;
	16'heee : data <= 32'h6384d101;
	16'heef : data <= 32'h6f309069;
	16'hef0 : data <= 32'hb700ff00;
	16'hef1 : data <= 32'h9380f00f;
	16'hef2 : data <= 32'h93e1f070;
	16'hef3 : data <= 32'hb70eff00;
	16'hef4 : data <= 32'h938efe7f;
	16'hef5 : data <= 32'h130ed016;
	16'hef6 : data <= 32'h6384d101;
	16'hef7 : data <= 32'h6f309067;
	16'hef8 : data <= 32'hb7f00ff0;
	16'hef9 : data <= 32'h9380f000;
	16'hefa : data <= 32'h93e1000f;
	16'hefb : data <= 32'hb7fe0ff0;
	16'hefc : data <= 32'h938efe0f;
	16'hefd : data <= 32'h130ee016;
	16'hefe : data <= 32'h6384d101;
	16'heff : data <= 32'h6f309065;
	16'hf00 : data <= 32'hb70001ff;
	16'hf01 : data <= 32'h938000f0;
	16'hf02 : data <= 32'h93e0000f;
	16'hf03 : data <= 32'hb70e01ff;
	16'hf04 : data <= 32'h938e0eff;
	16'hf05 : data <= 32'h130ef016;
	16'hf06 : data <= 32'h6384d001;
	16'hf07 : data <= 32'h6f309063;
	16'hf08 : data <= 32'h13020000;
	16'hf09 : data <= 32'hb710f00f;
	16'hf0a : data <= 32'h938000ff;
	16'hf0b : data <= 32'h93e1000f;
	16'hf0c : data <= 32'h13830100;
	16'hf0d : data <= 32'h13021200;
	16'hf0e : data <= 32'h93022000;
	16'hf0f : data <= 32'he31452fe;
	16'hf10 : data <= 32'hb71ef00f;
	16'hf11 : data <= 32'h938e0eff;
	16'hf12 : data <= 32'h130e0017;
	16'hf13 : data <= 32'h6304d301;
	16'hf14 : data <= 32'h6f305060;
	16'hf15 : data <= 32'h13020000;
	16'hf16 : data <= 32'hb700ff00;
	16'hf17 : data <= 32'h9380f00f;
	16'hf18 : data <= 32'h93e1f070;
	16'hf19 : data <= 32'h13000000;
	16'hf1a : data <= 32'h13830100;
	16'hf1b : data <= 32'h13021200;
	16'hf1c : data <= 32'h93022000;
	16'hf1d : data <= 32'he31252fe;
	16'hf1e : data <= 32'hb70eff00;
	16'hf1f : data <= 32'h938efe7f;
	16'hf20 : data <= 32'h130e1017;
	16'hf21 : data <= 32'h6304d301;
	16'hf22 : data <= 32'h6f30d05c;
	16'hf23 : data <= 32'h13020000;
	16'hf24 : data <= 32'hb7f00ff0;
	16'hf25 : data <= 32'h9380f000;
	16'hf26 : data <= 32'h93e1000f;
	16'hf27 : data <= 32'h13000000;
	16'hf28 : data <= 32'h13000000;
	16'hf29 : data <= 32'h13830100;
	16'hf2a : data <= 32'h13021200;
	16'hf2b : data <= 32'h93022000;
	16'hf2c : data <= 32'he31052fe;
	16'hf2d : data <= 32'hb7fe0ff0;
	16'hf2e : data <= 32'h938efe0f;
	16'hf2f : data <= 32'h130e2017;
	16'hf30 : data <= 32'h6304d301;
	16'hf31 : data <= 32'h6f301059;
	16'hf32 : data <= 32'h13020000;
	16'hf33 : data <= 32'hb710f00f;
	16'hf34 : data <= 32'h938000ff;
	16'hf35 : data <= 32'h93e1000f;
	16'hf36 : data <= 32'h13021200;
	16'hf37 : data <= 32'h93022000;
	16'hf38 : data <= 32'he31652fe;
	16'hf39 : data <= 32'hb71ef00f;
	16'hf3a : data <= 32'h938e0eff;
	16'hf3b : data <= 32'h130e3017;
	16'hf3c : data <= 32'h6384d101;
	16'hf3d : data <= 32'h6f301056;
	16'hf3e : data <= 32'h13020000;
	16'hf3f : data <= 32'hb700ff00;
	16'hf40 : data <= 32'h9380f00f;
	16'hf41 : data <= 32'h13000000;
	16'hf42 : data <= 32'h93e1f0f0;
	16'hf43 : data <= 32'h13021200;
	16'hf44 : data <= 32'h93022000;
	16'hf45 : data <= 32'he31452fe;
	16'hf46 : data <= 32'h930ef0ff;
	16'hf47 : data <= 32'h130e4017;
	16'hf48 : data <= 32'h6384d101;
	16'hf49 : data <= 32'h6f301053;
	16'hf4a : data <= 32'h13020000;
	16'hf4b : data <= 32'hb7f00ff0;
	16'hf4c : data <= 32'h9380f000;
	16'hf4d : data <= 32'h13000000;
	16'hf4e : data <= 32'h13000000;
	16'hf4f : data <= 32'h93e1000f;
	16'hf50 : data <= 32'h13021200;
	16'hf51 : data <= 32'h93022000;
	16'hf52 : data <= 32'he31252fe;
	16'hf53 : data <= 32'hb7fe0ff0;
	16'hf54 : data <= 32'h938efe0f;
	16'hf55 : data <= 32'h130e5017;
	16'hf56 : data <= 32'h6384d101;
	16'hf57 : data <= 32'h6f30904f;
	16'hf58 : data <= 32'h9360000f;
	16'hf59 : data <= 32'h930e000f;
	16'hf5a : data <= 32'h130e6017;
	16'hf5b : data <= 32'h6384d001;
	16'hf5c : data <= 32'h6f30504e;
	16'hf5d : data <= 32'hb700ff00;
	16'hf5e : data <= 32'h9380f00f;
	16'hf5f : data <= 32'h13e0f070;
	16'hf60 : data <= 32'h930e0000;
	16'hf61 : data <= 32'h130e7017;
	16'hf62 : data <= 32'h6304d001;
	16'hf63 : data <= 32'h6f30904c;
	16'hf64 : data <= 32'h97400000;
	16'hf65 : data <= 32'h93808029;
	16'hf66 : data <= 32'h1301a0fa;
	16'hf67 : data <= 32'h23802000;
	16'hf68 : data <= 32'h83810000;
	16'hf69 : data <= 32'h930ea0fa;
	16'hf6a : data <= 32'h130e8017;
	16'hf6b : data <= 32'h6384d101;
	16'hf6c : data <= 32'h6f30504a;
	16'hf6d : data <= 32'h97400000;
	16'hf6e : data <= 32'h93804027;
	16'hf6f : data <= 32'h13010000;
	16'hf70 : data <= 32'ha3802000;
	16'hf71 : data <= 32'h83811000;
	16'hf72 : data <= 32'h930e0000;
	16'hf73 : data <= 32'h130e9017;
	16'hf74 : data <= 32'h6384d101;
	16'hf75 : data <= 32'h6f301048;
	16'hf76 : data <= 32'h97400000;
	16'hf77 : data <= 32'h93800025;
	16'hf78 : data <= 32'h37f1ffff;
	16'hf79 : data <= 32'h130101fa;
	16'hf7a : data <= 32'h23812000;
	16'hf7b : data <= 32'h83912000;
	16'hf7c : data <= 32'hb7feffff;
	16'hf7d : data <= 32'h938e0efa;
	16'hf7e : data <= 32'h130ea017;
	16'hf7f : data <= 32'h6384d101;
	16'hf80 : data <= 32'h6f305045;
	16'hf81 : data <= 32'h97400000;
	16'hf82 : data <= 32'h93804022;
	16'hf83 : data <= 32'h1301a000;
	16'hf84 : data <= 32'ha3812000;
	16'hf85 : data <= 32'h83813000;
	16'hf86 : data <= 32'h930ea000;
	16'hf87 : data <= 32'h130ec017;
	16'hf88 : data <= 32'h6384d101;
	16'hf89 : data <= 32'h6f301043;
	16'hf8a : data <= 32'h97400000;
	16'hf8b : data <= 32'h93807020;
	16'hf8c : data <= 32'h1301a0fa;
	16'hf8d : data <= 32'ha38e20fe;
	16'hf8e : data <= 32'h8381d0ff;
	16'hf8f : data <= 32'h930ea0fa;
	16'hf90 : data <= 32'h130ed017;
	16'hf91 : data <= 32'h6384d101;
	16'hf92 : data <= 32'h6f30d040;
	16'hf93 : data <= 32'h97400000;
	16'hf94 : data <= 32'h9380301e;
	16'hf95 : data <= 32'h13010000;
	16'hf96 : data <= 32'h238f20fe;
	16'hf97 : data <= 32'h8381e0ff;
	16'hf98 : data <= 32'h930e0000;
	16'hf99 : data <= 32'h130ee017;
	16'hf9a : data <= 32'h6384d101;
	16'hf9b : data <= 32'h6f30903e;
	16'hf9c : data <= 32'h97400000;
	16'hf9d : data <= 32'h9380f01b;
	16'hf9e : data <= 32'h130100fa;
	16'hf9f : data <= 32'ha38f20fe;
	16'hfa0 : data <= 32'h8381f0ff;
	16'hfa1 : data <= 32'h930e00fa;
	16'hfa2 : data <= 32'h130ef017;
	16'hfa3 : data <= 32'h6384d101;
	16'hfa4 : data <= 32'h6f30503c;
	16'hfa5 : data <= 32'h97400000;
	16'hfa6 : data <= 32'h9380b019;
	16'hfa7 : data <= 32'h1301a000;
	16'hfa8 : data <= 32'h23802000;
	16'hfa9 : data <= 32'h83810000;
	16'hfaa : data <= 32'h930ea000;
	16'hfab : data <= 32'h130e0018;
	16'hfac : data <= 32'h6384d101;
	16'hfad : data <= 32'h6f30103a;
	16'hfae : data <= 32'h97400000;
	16'hfaf : data <= 32'h93808017;
	16'hfb0 : data <= 32'h37513412;
	16'hfb1 : data <= 32'h13018167;
	16'hfb2 : data <= 32'h138200fe;
	16'hfb3 : data <= 32'h23002202;
	16'hfb4 : data <= 32'h83810000;
	16'hfb5 : data <= 32'h930e8007;
	16'hfb6 : data <= 32'h130e1018;
	16'hfb7 : data <= 32'h6384d101;
	16'hfb8 : data <= 32'h6f305037;
	16'hfb9 : data <= 32'h97400000;
	16'hfba : data <= 32'h9380c014;
	16'hfbb : data <= 32'h37310000;
	16'hfbc : data <= 32'h13018109;
	16'hfbd : data <= 32'h9380a0ff;
	16'hfbe : data <= 32'ha3832000;
	16'hfbf : data <= 32'h17420000;
	16'hfc0 : data <= 32'h13025213;
	16'hfc1 : data <= 32'h83010200;
	16'hfc2 : data <= 32'h930e80f9;
	16'hfc3 : data <= 32'h130e2018;
	16'hfc4 : data <= 32'h6384d101;
	16'hfc5 : data <= 32'h6f301034;
	16'hfc6 : data <= 32'h130e3018;
	16'hfc7 : data <= 32'h13020000;
	16'hfc8 : data <= 32'h9300d0fd;
	16'hfc9 : data <= 32'h17410000;
	16'hfca : data <= 32'h13014110;
	16'hfcb : data <= 32'h23001100;
	16'hfcc : data <= 32'h83010100;
	16'hfcd : data <= 32'h930ed0fd;
	16'hfce : data <= 32'h6384d101;
	16'hfcf : data <= 32'h6f309031;
	16'hfd0 : data <= 32'h13021200;
	16'hfd1 : data <= 32'h93022000;
	16'hfd2 : data <= 32'he31c52fc;
	16'hfd3 : data <= 32'h130e4018;
	16'hfd4 : data <= 32'h13020000;
	16'hfd5 : data <= 32'h9300d0fc;
	16'hfd6 : data <= 32'h17410000;
	16'hfd7 : data <= 32'h1301010d;
	16'hfd8 : data <= 32'h13000000;
	16'hfd9 : data <= 32'ha3001100;
	16'hfda : data <= 32'h83011100;
	16'hfdb : data <= 32'h930ed0fc;
	16'hfdc : data <= 32'h6384d101;
	16'hfdd : data <= 32'h6f30102e;
	16'hfde : data <= 32'h13021200;
	16'hfdf : data <= 32'h93022000;
	16'hfe0 : data <= 32'he31a52fc;
	16'hfe1 : data <= 32'h130e5018;
	16'hfe2 : data <= 32'h13020000;
	16'hfe3 : data <= 32'h9300c0fc;
	16'hfe4 : data <= 32'h17410000;
	16'hfe5 : data <= 32'h13018109;
	16'hfe6 : data <= 32'h13000000;
	16'hfe7 : data <= 32'h13000000;
	16'hfe8 : data <= 32'h23011100;
	16'hfe9 : data <= 32'h83012100;
	16'hfea : data <= 32'h930ec0fc;
	16'hfeb : data <= 32'h6384d101;
	16'hfec : data <= 32'h6f30502a;
	16'hfed : data <= 32'h13021200;
	16'hfee : data <= 32'h93022000;
	16'hfef : data <= 32'he31852fc;
	16'hff0 : data <= 32'h130e6018;
	16'hff1 : data <= 32'h13020000;
	16'hff2 : data <= 32'h9300c0fb;
	16'hff3 : data <= 32'h13000000;
	16'hff4 : data <= 32'h17410000;
	16'hff5 : data <= 32'h13018105;
	16'hff6 : data <= 32'ha3011100;
	16'hff7 : data <= 32'h83013100;
	16'hff8 : data <= 32'h930ec0fb;
	16'hff9 : data <= 32'h6384d101;
	16'hffa : data <= 32'h6f30d026;
	16'hffb : data <= 32'h13021200;
	16'hffc : data <= 32'h93022000;
	16'hffd : data <= 32'he31a52fc;
	16'hffe : data <= 32'h130e7018;
	16'hfff : data <= 32'h13020000;
	16'h1000 : data <= 32'h9300b0fb;
	16'h1001 : data <= 32'h13000000;
	16'h1002 : data <= 32'h17410000;
	16'h1003 : data <= 32'h13010102;
	16'h1004 : data <= 32'h13000000;
	16'h1005 : data <= 32'h23021100;
	16'h1006 : data <= 32'h83014100;
	16'h1007 : data <= 32'h930eb0fb;
	16'h1008 : data <= 32'h6384d101;
	16'h1009 : data <= 32'h6f301023;
	16'h100a : data <= 32'h13021200;
	16'h100b : data <= 32'h93022000;
	16'h100c : data <= 32'he31852fc;
	16'h100d : data <= 32'h130e8018;
	16'h100e : data <= 32'h13020000;
	16'h100f : data <= 32'h9300b0fa;
	16'h1010 : data <= 32'h13000000;
	16'h1011 : data <= 32'h13000000;
	16'h1012 : data <= 32'h17410000;
	16'h1013 : data <= 32'h130101fe;
	16'h1014 : data <= 32'ha3021100;
	16'h1015 : data <= 32'h83015100;
	16'h1016 : data <= 32'h930eb0fa;
	16'h1017 : data <= 32'h6384d101;
	16'h1018 : data <= 32'h6f30501f;
	16'h1019 : data <= 32'h13021200;
	16'h101a : data <= 32'h93022000;
	16'h101b : data <= 32'he31852fc;
	16'h101c : data <= 32'h130e9018;
	16'h101d : data <= 32'h13020000;
	16'h101e : data <= 32'h17410000;
	16'h101f : data <= 32'h130101fb;
	16'h1020 : data <= 32'h93003003;
	16'h1021 : data <= 32'h23001100;
	16'h1022 : data <= 32'h83010100;
	16'h1023 : data <= 32'h930e3003;
	16'h1024 : data <= 32'h6384d101;
	16'h1025 : data <= 32'h6f30101c;
	16'h1026 : data <= 32'h13021200;
	16'h1027 : data <= 32'h93022000;
	16'h1028 : data <= 32'he31c52fc;
	16'h1029 : data <= 32'h130ea018;
	16'h102a : data <= 32'h13020000;
	16'h102b : data <= 32'h17410000;
	16'h102c : data <= 32'h1301c1f7;
	16'h102d : data <= 32'h93003002;
	16'h102e : data <= 32'h13000000;
	16'h102f : data <= 32'ha3001100;
	16'h1030 : data <= 32'h83011100;
	16'h1031 : data <= 32'h930e3002;
	16'h1032 : data <= 32'h6384d101;
	16'h1033 : data <= 32'h6f309018;
	16'h1034 : data <= 32'h13021200;
	16'h1035 : data <= 32'h93022000;
	16'h1036 : data <= 32'he31a52fc;
	16'h1037 : data <= 32'h130eb018;
	16'h1038 : data <= 32'h13020000;
	16'h1039 : data <= 32'h17410000;
	16'h103a : data <= 32'h130141f4;
	16'h103b : data <= 32'h93002002;
	16'h103c : data <= 32'h13000000;
	16'h103d : data <= 32'h13000000;
	16'h103e : data <= 32'h23011100;
	16'h103f : data <= 32'h83012100;
	16'h1040 : data <= 32'h930e2002;
	16'h1041 : data <= 32'h6384d101;
	16'h1042 : data <= 32'h6f30d014;
	16'h1043 : data <= 32'h13021200;
	16'h1044 : data <= 32'h93022000;
	16'h1045 : data <= 32'he31852fc;
	16'h1046 : data <= 32'h130ec018;
	16'h1047 : data <= 32'h13020000;
	16'h1048 : data <= 32'h17410000;
	16'h1049 : data <= 32'h130181f0;
	16'h104a : data <= 32'h13000000;
	16'h104b : data <= 32'h93002001;
	16'h104c : data <= 32'ha3011100;
	16'h104d : data <= 32'h83013100;
	16'h104e : data <= 32'h930e2001;
	16'h104f : data <= 32'h6384d101;
	16'h1050 : data <= 32'h6f305011;
	16'h1051 : data <= 32'h13021200;
	16'h1052 : data <= 32'h93022000;
	16'h1053 : data <= 32'he31a52fc;
	16'h1054 : data <= 32'h130ed018;
	16'h1055 : data <= 32'h13020000;
	16'h1056 : data <= 32'h17410000;
	16'h1057 : data <= 32'h130101ed;
	16'h1058 : data <= 32'h13000000;
	16'h1059 : data <= 32'h93001001;
	16'h105a : data <= 32'h13000000;
	16'h105b : data <= 32'h23021100;
	16'h105c : data <= 32'h83014100;
	16'h105d : data <= 32'h930e1001;
	16'h105e : data <= 32'h6384d101;
	16'h105f : data <= 32'h6f30900d;
	16'h1060 : data <= 32'h13021200;
	16'h1061 : data <= 32'h93022000;
	16'h1062 : data <= 32'he31852fc;
	16'h1063 : data <= 32'h130ee018;
	16'h1064 : data <= 32'h13020000;
	16'h1065 : data <= 32'h17410000;
	16'h1066 : data <= 32'h130141e9;
	16'h1067 : data <= 32'h13000000;
	16'h1068 : data <= 32'h13000000;
	16'h1069 : data <= 32'h93001000;
	16'h106a : data <= 32'ha3021100;
	16'h106b : data <= 32'h83015100;
	16'h106c : data <= 32'h930e1000;
	16'h106d : data <= 32'h6384d101;
	16'h106e : data <= 32'h6f30d009;
	16'h106f : data <= 32'h13021200;
	16'h1070 : data <= 32'h93022000;
	16'h1071 : data <= 32'he31852fc;
	16'h1072 : data <= 32'h1305f00e;
	16'h1073 : data <= 32'h97450000;
	16'h1074 : data <= 32'h9385c5e5;
	16'h1075 : data <= 32'ha381a500;
	16'h1076 : data <= 32'h97400000;
	16'h1077 : data <= 32'h9380a0e5;
	16'h1078 : data <= 32'h1301a00a;
	16'h1079 : data <= 32'h23902000;
	16'h107a : data <= 32'h83910000;
	16'h107b : data <= 32'h930ea00a;
	16'h107c : data <= 32'h130ef018;
	16'h107d : data <= 32'h6384d101;
	16'h107e : data <= 32'h6f30d005;
	16'h107f : data <= 32'h97400000;
	16'h1080 : data <= 32'h938060e3;
	16'h1081 : data <= 32'h37b1ffff;
	16'h1082 : data <= 32'h130101a0;
	16'h1083 : data <= 32'h23912000;
	16'h1084 : data <= 32'h83912000;
	16'h1085 : data <= 32'hb7beffff;
	16'h1086 : data <= 32'h938e0ea0;
	16'h1087 : data <= 32'h130e0019;
	16'h1088 : data <= 32'h6384d101;
	16'h1089 : data <= 32'h6f301003;
	16'h108a : data <= 32'h97400000;
	16'h108b : data <= 32'h9380a0e0;
	16'h108c : data <= 32'h3711efbe;
	16'h108d : data <= 32'h130101aa;
	16'h108e : data <= 32'h23922000;
	16'h108f : data <= 32'h83a14000;
	16'h1090 : data <= 32'hb71eefbe;
	16'h1091 : data <= 32'h938e0eaa;
	16'h1092 : data <= 32'h130e1019;
	16'h1093 : data <= 32'h6384d101;
	16'h1094 : data <= 32'h6f305000;
	16'h1095 : data <= 32'h97400000;
	16'h1096 : data <= 32'h9380e0dd;
	16'h1097 : data <= 32'h37a1ffff;
	16'h1098 : data <= 32'h1301a100;
	16'h1099 : data <= 32'h23932000;
	16'h109a : data <= 32'h83916000;
	16'h109b : data <= 32'hb7aeffff;
	16'h109c : data <= 32'h938eae00;
	16'h109d : data <= 32'h130e2019;
	16'h109e : data <= 32'h6384d101;
	16'h109f : data <= 32'h6f30807d;
	16'h10a0 : data <= 32'h97400000;
	16'h10a1 : data <= 32'h938000dc;
	16'h10a2 : data <= 32'h1301a00a;
	16'h10a3 : data <= 32'h239d20fe;
	16'h10a4 : data <= 32'h8391a0ff;
	16'h10a5 : data <= 32'h930ea00a;
	16'h10a6 : data <= 32'h130e3019;
	16'h10a7 : data <= 32'h6384d101;
	16'h10a8 : data <= 32'h6f30407b;
	16'h10a9 : data <= 32'h97400000;
	16'h10aa : data <= 32'h9380c0d9;
	16'h10ab : data <= 32'h37b1ffff;
	16'h10ac : data <= 32'h130101a0;
	16'h10ad : data <= 32'h239e20fe;
	16'h10ae : data <= 32'h8391c0ff;
	16'h10af : data <= 32'hb7beffff;
	16'h10b0 : data <= 32'h938e0ea0;
	16'h10b1 : data <= 32'h130e4019;
	16'h10b2 : data <= 32'h6384d101;
	16'h10b3 : data <= 32'h6f308078;
	16'h10b4 : data <= 32'h97400000;
	16'h10b5 : data <= 32'h938000d7;
	16'h10b6 : data <= 32'h37110000;
	16'h10b7 : data <= 32'h130101aa;
	16'h10b8 : data <= 32'h239f20fe;
	16'h10b9 : data <= 32'h8391e0ff;
	16'h10ba : data <= 32'hb71e0000;
	16'h10bb : data <= 32'h938e0eaa;
	16'h10bc : data <= 32'h130e5019;
	16'h10bd : data <= 32'h6384d101;
	16'h10be : data <= 32'h6f30c075;
	16'h10bf : data <= 32'h97400000;
	16'h10c0 : data <= 32'h938040d4;
	16'h10c1 : data <= 32'h37a1ffff;
	16'h10c2 : data <= 32'h1301a100;
	16'h10c3 : data <= 32'h23902000;
	16'h10c4 : data <= 32'h83910000;
	16'h10c5 : data <= 32'hb7aeffff;
	16'h10c6 : data <= 32'h938eae00;
	16'h10c7 : data <= 32'h130e6019;
	16'h10c8 : data <= 32'h6384d101;
	16'h10c9 : data <= 32'h6f300073;
	16'h10ca : data <= 32'h97400000;
	16'h10cb : data <= 32'h9380a0d1;
	16'h10cc : data <= 32'h37513412;
	16'h10cd : data <= 32'h13018167;
	16'h10ce : data <= 32'h138200fe;
	16'h10cf : data <= 32'h23102202;
	16'h10d0 : data <= 32'h83910000;
	16'h10d1 : data <= 32'hb75e0000;
	16'h10d2 : data <= 32'h938e8e67;
	16'h10d3 : data <= 32'h130e7019;
	16'h10d4 : data <= 32'h6384d101;
	16'h10d5 : data <= 32'h6f300070;
	16'h10d6 : data <= 32'h97400000;
	16'h10d7 : data <= 32'h9380a0ce;
	16'h10d8 : data <= 32'h37310000;
	16'h10d9 : data <= 32'h13018109;
	16'h10da : data <= 32'h9380b0ff;
	16'h10db : data <= 32'ha3932000;
	16'h10dc : data <= 32'h17420000;
	16'h10dd : data <= 32'h130242cd;
	16'h10de : data <= 32'h83110200;
	16'h10df : data <= 32'hb73e0000;
	16'h10e0 : data <= 32'h938e8e09;
	16'h10e1 : data <= 32'h130e8019;
	16'h10e2 : data <= 32'h6384d101;
	16'h10e3 : data <= 32'h6f30806c;
	16'h10e4 : data <= 32'h130e9019;
	16'h10e5 : data <= 32'h13020000;
	16'h10e6 : data <= 32'hb7d0ffff;
	16'h10e7 : data <= 32'h9380d0cd;
	16'h10e8 : data <= 32'h17410000;
	16'h10e9 : data <= 32'h130121c9;
	16'h10ea : data <= 32'h23101100;
	16'h10eb : data <= 32'h83110100;
	16'h10ec : data <= 32'hb7deffff;
	16'h10ed : data <= 32'h938edecd;
	16'h10ee : data <= 32'h6384d101;
	16'h10ef : data <= 32'h6f308069;
	16'h10f0 : data <= 32'h13021200;
	16'h10f1 : data <= 32'h93022000;
	16'h10f2 : data <= 32'he31852fc;
	16'h10f3 : data <= 32'h130ea019;
	16'h10f4 : data <= 32'h13020000;
	16'h10f5 : data <= 32'hb7c0ffff;
	16'h10f6 : data <= 32'h9380d0cc;
	16'h10f7 : data <= 32'h17410000;
	16'h10f8 : data <= 32'h130161c5;
	16'h10f9 : data <= 32'h13000000;
	16'h10fa : data <= 32'h23111100;
	16'h10fb : data <= 32'h83112100;
	16'h10fc : data <= 32'hb7ceffff;
	16'h10fd : data <= 32'h938edecc;
	16'h10fe : data <= 32'h6384d101;
	16'h10ff : data <= 32'h6f308065;
	16'h1100 : data <= 32'h13021200;
	16'h1101 : data <= 32'h93022000;
	16'h1102 : data <= 32'he31652fc;
	16'h1103 : data <= 32'h130eb019;
	16'h1104 : data <= 32'h13020000;
	16'h1105 : data <= 32'hb7c0ffff;
	16'h1106 : data <= 32'h9380c0bc;
	16'h1107 : data <= 32'h17410000;
	16'h1108 : data <= 32'h130161c1;
	16'h1109 : data <= 32'h13000000;
	16'h110a : data <= 32'h13000000;
	16'h110b : data <= 32'h23121100;
	16'h110c : data <= 32'h83114100;
	16'h110d : data <= 32'hb7ceffff;
	16'h110e : data <= 32'h938ecebc;
	16'h110f : data <= 32'h6384d101;
	16'h1110 : data <= 32'h6f304061;
	16'h1111 : data <= 32'h13021200;
	16'h1112 : data <= 32'h93022000;
	16'h1113 : data <= 32'he31452fc;
	16'h1114 : data <= 32'h130ec019;
	16'h1115 : data <= 32'h13020000;
	16'h1116 : data <= 32'hb7b0ffff;
	16'h1117 : data <= 32'h9380c0bb;
	16'h1118 : data <= 32'h13000000;
	16'h1119 : data <= 32'h17410000;
	16'h111a : data <= 32'h1301e1bc;
	16'h111b : data <= 32'h23131100;
	16'h111c : data <= 32'h83116100;
	16'h111d : data <= 32'hb7beffff;
	16'h111e : data <= 32'h938ecebb;
	16'h111f : data <= 32'h6384d101;
	16'h1120 : data <= 32'h6f30405d;
	16'h1121 : data <= 32'h13021200;
	16'h1122 : data <= 32'h93022000;
	16'h1123 : data <= 32'he31652fc;
	16'h1124 : data <= 32'h130ed019;
	16'h1125 : data <= 32'h13020000;
	16'h1126 : data <= 32'hb7b0ffff;
	16'h1127 : data <= 32'h9380b0ab;
	16'h1128 : data <= 32'h13000000;
	16'h1129 : data <= 32'h17410000;
	16'h112a : data <= 32'h1301e1b8;
	16'h112b : data <= 32'h13000000;
	16'h112c : data <= 32'h23141100;
	16'h112d : data <= 32'h83118100;
	16'h112e : data <= 32'hb7beffff;
	16'h112f : data <= 32'h938ebeab;
	16'h1130 : data <= 32'h6384d101;
	16'h1131 : data <= 32'h6f300059;
	16'h1132 : data <= 32'h13021200;
	16'h1133 : data <= 32'h93022000;
	16'h1134 : data <= 32'he31452fc;
	16'h1135 : data <= 32'h130ee019;
	16'h1136 : data <= 32'h13020000;
	16'h1137 : data <= 32'hb7e0ffff;
	16'h1138 : data <= 32'h9380b0aa;
	16'h1139 : data <= 32'h13000000;
	16'h113a : data <= 32'h13000000;
	16'h113b : data <= 32'h17410000;
	16'h113c : data <= 32'h130161b4;
	16'h113d : data <= 32'h23151100;
	16'h113e : data <= 32'h8311a100;
	16'h113f : data <= 32'hb7eeffff;
	16'h1140 : data <= 32'h938ebeaa;
	16'h1141 : data <= 32'h6384d101;
	16'h1142 : data <= 32'h6f30c054;
	16'h1143 : data <= 32'h13021200;
	16'h1144 : data <= 32'h93022000;
	16'h1145 : data <= 32'he31452fc;
	16'h1146 : data <= 32'h130ef019;
	16'h1147 : data <= 32'h13020000;
	16'h1148 : data <= 32'h17410000;
	16'h1149 : data <= 32'h130121b1;
	16'h114a : data <= 32'hb7200000;
	16'h114b : data <= 32'h93803023;
	16'h114c : data <= 32'h23101100;
	16'h114d : data <= 32'h83110100;
	16'h114e : data <= 32'hb72e0000;
	16'h114f : data <= 32'h938e3e23;
	16'h1150 : data <= 32'h6384d101;
	16'h1151 : data <= 32'h6f300051;
	16'h1152 : data <= 32'h13021200;
	16'h1153 : data <= 32'h93022000;
	16'h1154 : data <= 32'he31852fc;
	16'h1155 : data <= 32'h130e001a;
	16'h1156 : data <= 32'h13020000;
	16'h1157 : data <= 32'h17410000;
	16'h1158 : data <= 32'h130161ad;
	16'h1159 : data <= 32'hb7100000;
	16'h115a : data <= 32'h93803022;
	16'h115b : data <= 32'h13000000;
	16'h115c : data <= 32'h23111100;
	16'h115d : data <= 32'h83112100;
	16'h115e : data <= 32'hb71e0000;
	16'h115f : data <= 32'h938e3e22;
	16'h1160 : data <= 32'h6384d101;
	16'h1161 : data <= 32'h6f30004d;
	16'h1162 : data <= 32'h13021200;
	16'h1163 : data <= 32'h93022000;
	16'h1164 : data <= 32'he31652fc;
	16'h1165 : data <= 32'h130e101a;
	16'h1166 : data <= 32'h13020000;
	16'h1167 : data <= 32'h17410000;
	16'h1168 : data <= 32'h130161a9;
	16'h1169 : data <= 32'hb7100000;
	16'h116a : data <= 32'h93802012;
	16'h116b : data <= 32'h13000000;
	16'h116c : data <= 32'h13000000;
	16'h116d : data <= 32'h23121100;
	16'h116e : data <= 32'h83114100;
	16'h116f : data <= 32'hb71e0000;
	16'h1170 : data <= 32'h938e2e12;
	16'h1171 : data <= 32'h6384d101;
	16'h1172 : data <= 32'h6f30c048;
	16'h1173 : data <= 32'h13021200;
	16'h1174 : data <= 32'h93022000;
	16'h1175 : data <= 32'he31452fc;
	16'h1176 : data <= 32'h130e201a;
	16'h1177 : data <= 32'h13020000;
	16'h1178 : data <= 32'h17410000;
	16'h1179 : data <= 32'h130121a5;
	16'h117a : data <= 32'h13000000;
	16'h117b : data <= 32'h93002011;
	16'h117c : data <= 32'h23131100;
	16'h117d : data <= 32'h83116100;
	16'h117e : data <= 32'h930e2011;
	16'h117f : data <= 32'h6384d101;
	16'h1180 : data <= 32'h6f304045;
	16'h1181 : data <= 32'h13021200;
	16'h1182 : data <= 32'h93022000;
	16'h1183 : data <= 32'he31a52fc;
	16'h1184 : data <= 32'h130e301a;
	16'h1185 : data <= 32'h13020000;
	16'h1186 : data <= 32'h17410000;
	16'h1187 : data <= 32'h1301a1a1;
	16'h1188 : data <= 32'h13000000;
	16'h1189 : data <= 32'h93001001;
	16'h118a : data <= 32'h13000000;
	16'h118b : data <= 32'h23141100;
	16'h118c : data <= 32'h83118100;
	16'h118d : data <= 32'h930e1001;
	16'h118e : data <= 32'h6384d101;
	16'h118f : data <= 32'h6f308041;
	16'h1190 : data <= 32'h13021200;
	16'h1191 : data <= 32'h93022000;
	16'h1192 : data <= 32'he31852fc;
	16'h1193 : data <= 32'h130e401a;
	16'h1194 : data <= 32'h13020000;
	16'h1195 : data <= 32'h17410000;
	16'h1196 : data <= 32'h1301e19d;
	16'h1197 : data <= 32'h13000000;
	16'h1198 : data <= 32'h13000000;
	16'h1199 : data <= 32'hb7300000;
	16'h119a : data <= 32'h93801000;
	16'h119b : data <= 32'h23151100;
	16'h119c : data <= 32'h8311a100;
	16'h119d : data <= 32'hb73e0000;
	16'h119e : data <= 32'h938e1e00;
	16'h119f : data <= 32'h6384d101;
	16'h11a0 : data <= 32'h6f30403d;
	16'h11a1 : data <= 32'h13021200;
	16'h11a2 : data <= 32'h93022000;
	16'h11a3 : data <= 32'he31452fc;
	16'h11a4 : data <= 32'h37c50000;
	16'h11a5 : data <= 32'h1305f5ee;
	16'h11a6 : data <= 32'h97450000;
	16'h11a7 : data <= 32'h9385a599;
	16'h11a8 : data <= 32'h2393a500;
	16'h11a9 : data <= 32'h93001000;
	16'h11aa : data <= 32'h13010000;
	16'h11ab : data <= 32'hb3912000;
	16'h11ac : data <= 32'h930e1000;
	16'h11ad : data <= 32'h130e501a;
	16'h11ae : data <= 32'h6384d101;
	16'h11af : data <= 32'h6f308039;
	16'h11b0 : data <= 32'h93001000;
	16'h11b1 : data <= 32'h13011000;
	16'h11b2 : data <= 32'hb3912000;
	16'h11b3 : data <= 32'h930e2000;
	16'h11b4 : data <= 32'h130e601a;
	16'h11b5 : data <= 32'h6384d101;
	16'h11b6 : data <= 32'h6f30c037;
	16'h11b7 : data <= 32'h93001000;
	16'h11b8 : data <= 32'h13017000;
	16'h11b9 : data <= 32'hb3912000;
	16'h11ba : data <= 32'h930e0008;
	16'h11bb : data <= 32'h130e701a;
	16'h11bc : data <= 32'h6384d101;
	16'h11bd : data <= 32'h6f300036;
	16'h11be : data <= 32'h93001000;
	16'h11bf : data <= 32'h1301e000;
	16'h11c0 : data <= 32'hb3912000;
	16'h11c1 : data <= 32'hb74e0000;
	16'h11c2 : data <= 32'h130e801a;
	16'h11c3 : data <= 32'h6384d101;
	16'h11c4 : data <= 32'h6f304034;
	16'h11c5 : data <= 32'h93001000;
	16'h11c6 : data <= 32'h1301f001;
	16'h11c7 : data <= 32'hb3912000;
	16'h11c8 : data <= 32'hb70e0080;
	16'h11c9 : data <= 32'h130e901a;
	16'h11ca : data <= 32'h6384d101;
	16'h11cb : data <= 32'h6f308032;
	16'h11cc : data <= 32'h9300f0ff;
	16'h11cd : data <= 32'h13010000;
	16'h11ce : data <= 32'hb3912000;
	16'h11cf : data <= 32'h930ef0ff;
	16'h11d0 : data <= 32'h130ea01a;
	16'h11d1 : data <= 32'h6384d101;
	16'h11d2 : data <= 32'h6f30c030;
	16'h11d3 : data <= 32'h9300f0ff;
	16'h11d4 : data <= 32'h13011000;
	16'h11d5 : data <= 32'hb3912000;
	16'h11d6 : data <= 32'h930ee0ff;
	16'h11d7 : data <= 32'h130eb01a;
	16'h11d8 : data <= 32'h6384d101;
	16'h11d9 : data <= 32'h6f30002f;
	16'h11da : data <= 32'h9300f0ff;
	16'h11db : data <= 32'h13017000;
	16'h11dc : data <= 32'hb3912000;
	16'h11dd : data <= 32'h930e00f8;
	16'h11de : data <= 32'h130ec01a;
	16'h11df : data <= 32'h6384d101;
	16'h11e0 : data <= 32'h6f30402d;
	16'h11e1 : data <= 32'h9300f0ff;
	16'h11e2 : data <= 32'h1301e000;
	16'h11e3 : data <= 32'hb3912000;
	16'h11e4 : data <= 32'hb7ceffff;
	16'h11e5 : data <= 32'h130ed01a;
	16'h11e6 : data <= 32'h6384d101;
	16'h11e7 : data <= 32'h6f30802b;
	16'h11e8 : data <= 32'h9300f0ff;
	16'h11e9 : data <= 32'h1301f001;
	16'h11ea : data <= 32'hb3912000;
	16'h11eb : data <= 32'hb70e0080;
	16'h11ec : data <= 32'h130ee01a;
	16'h11ed : data <= 32'h6384d101;
	16'h11ee : data <= 32'h6f30c029;
	16'h11ef : data <= 32'hb7202121;
	16'h11f0 : data <= 32'h93801012;
	16'h11f1 : data <= 32'h13010000;
	16'h11f2 : data <= 32'hb3912000;
	16'h11f3 : data <= 32'hb72e2121;
	16'h11f4 : data <= 32'h938e1e12;
	16'h11f5 : data <= 32'h130ef01a;
	16'h11f6 : data <= 32'h6384d101;
	16'h11f7 : data <= 32'h6f308027;
	16'h11f8 : data <= 32'hb7202121;
	16'h11f9 : data <= 32'h93801012;
	16'h11fa : data <= 32'h13011000;
	16'h11fb : data <= 32'hb3912000;
	16'h11fc : data <= 32'hb74e4242;
	16'h11fd : data <= 32'h938e2e24;
	16'h11fe : data <= 32'h130e001b;
	16'h11ff : data <= 32'h6384d101;
	16'h1200 : data <= 32'h6f304025;
	16'h1201 : data <= 32'hb7202121;
	16'h1202 : data <= 32'h93801012;
	16'h1203 : data <= 32'h13017000;
	16'h1204 : data <= 32'hb3912000;
	16'h1205 : data <= 32'hb79e9090;
	16'h1206 : data <= 32'h938e0e08;
	16'h1207 : data <= 32'h130e101b;
	16'h1208 : data <= 32'h6384d101;
	16'h1209 : data <= 32'h6f300023;
	16'h120a : data <= 32'hb7202121;
	16'h120b : data <= 32'h93801012;
	16'h120c : data <= 32'h1301e000;
	16'h120d : data <= 32'hb3912000;
	16'h120e : data <= 32'hb74e4848;
	16'h120f : data <= 32'h130e201b;
	16'h1210 : data <= 32'h6384d101;
	16'h1211 : data <= 32'h6f300021;
	16'h1212 : data <= 32'hb7202121;
	16'h1213 : data <= 32'h93801012;
	16'h1214 : data <= 32'h1301f001;
	16'h1215 : data <= 32'hb3912000;
	16'h1216 : data <= 32'hb70e0080;
	16'h1217 : data <= 32'h130e301b;
	16'h1218 : data <= 32'h6384d101;
	16'h1219 : data <= 32'h6f30001f;
	16'h121a : data <= 32'hb7202121;
	16'h121b : data <= 32'h93801012;
	16'h121c : data <= 32'h130100fe;
	16'h121d : data <= 32'hb3912000;
	16'h121e : data <= 32'hb72e2121;
	16'h121f : data <= 32'h938e1e12;
	16'h1220 : data <= 32'h130e401b;
	16'h1221 : data <= 32'h6384d101;
	16'h1222 : data <= 32'h6f30c01c;
	16'h1223 : data <= 32'hb7202121;
	16'h1224 : data <= 32'h93801012;
	16'h1225 : data <= 32'h130110fe;
	16'h1226 : data <= 32'hb3912000;
	16'h1227 : data <= 32'hb74e4242;
	16'h1228 : data <= 32'h938e2e24;
	16'h1229 : data <= 32'h130e501b;
	16'h122a : data <= 32'h6384d101;
	16'h122b : data <= 32'h6f30801a;
	16'h122c : data <= 32'hb7202121;
	16'h122d : data <= 32'h93801012;
	16'h122e : data <= 32'h130170fe;
	16'h122f : data <= 32'hb3912000;
	16'h1230 : data <= 32'hb79e9090;
	16'h1231 : data <= 32'h938e0e08;
	16'h1232 : data <= 32'h130e601b;
	16'h1233 : data <= 32'h6384d101;
	16'h1234 : data <= 32'h6f304018;
	16'h1235 : data <= 32'hb7202121;
	16'h1236 : data <= 32'h93801012;
	16'h1237 : data <= 32'h1301e0fe;
	16'h1238 : data <= 32'hb3912000;
	16'h1239 : data <= 32'hb74e4848;
	16'h123a : data <= 32'h130e701b;
	16'h123b : data <= 32'h6384d101;
	16'h123c : data <= 32'h6f304016;
	16'h123d : data <= 32'hb7202121;
	16'h123e : data <= 32'h93800012;
	16'h123f : data <= 32'h1301f0ff;
	16'h1240 : data <= 32'hb3912000;
	16'h1241 : data <= 32'h930e0000;
	16'h1242 : data <= 32'h130e801b;
	16'h1243 : data <= 32'h6384d101;
	16'h1244 : data <= 32'h6f304014;
	16'h1245 : data <= 32'h93001000;
	16'h1246 : data <= 32'h13017000;
	16'h1247 : data <= 32'hb3902000;
	16'h1248 : data <= 32'h930e0008;
	16'h1249 : data <= 32'h130e901b;
	16'h124a : data <= 32'h6384d001;
	16'h124b : data <= 32'h6f308012;
	16'h124c : data <= 32'h93001000;
	16'h124d : data <= 32'h1301e000;
	16'h124e : data <= 32'h33912000;
	16'h124f : data <= 32'hb74e0000;
	16'h1250 : data <= 32'h130ea01b;
	16'h1251 : data <= 32'h6304d101;
	16'h1252 : data <= 32'h6f30c010;
	16'h1253 : data <= 32'h93003000;
	16'h1254 : data <= 32'hb3901000;
	16'h1255 : data <= 32'h930e8001;
	16'h1256 : data <= 32'h130eb01b;
	16'h1257 : data <= 32'h6384d001;
	16'h1258 : data <= 32'h6f30400f;
	16'h1259 : data <= 32'h13020000;
	16'h125a : data <= 32'h93001000;
	16'h125b : data <= 32'h13017000;
	16'h125c : data <= 32'hb3912000;
	16'h125d : data <= 32'h13830100;
	16'h125e : data <= 32'h13021200;
	16'h125f : data <= 32'h93022000;
	16'h1260 : data <= 32'he31452fe;
	16'h1261 : data <= 32'h930e0008;
	16'h1262 : data <= 32'h130ec01b;
	16'h1263 : data <= 32'h6304d301;
	16'h1264 : data <= 32'h6f30400c;
	16'h1265 : data <= 32'h13020000;
	16'h1266 : data <= 32'h93001000;
	16'h1267 : data <= 32'h1301e000;
	16'h1268 : data <= 32'hb3912000;
	16'h1269 : data <= 32'h13000000;
	16'h126a : data <= 32'h13830100;
	16'h126b : data <= 32'h13021200;
	16'h126c : data <= 32'h93022000;
	16'h126d : data <= 32'he31252fe;
	16'h126e : data <= 32'hb74e0000;
	16'h126f : data <= 32'h130ed01b;
	16'h1270 : data <= 32'h6304d301;
	16'h1271 : data <= 32'h6f300009;
	16'h1272 : data <= 32'h13020000;
	16'h1273 : data <= 32'h93001000;
	16'h1274 : data <= 32'h1301f001;
	16'h1275 : data <= 32'hb3912000;
	16'h1276 : data <= 32'h13000000;
	16'h1277 : data <= 32'h13000000;
	16'h1278 : data <= 32'h13830100;
	16'h1279 : data <= 32'h13021200;
	16'h127a : data <= 32'h93022000;
	16'h127b : data <= 32'he31052fe;
	16'h127c : data <= 32'hb70e0080;
	16'h127d : data <= 32'h130ee01b;
	16'h127e : data <= 32'h6304d301;
	16'h127f : data <= 32'h6f308005;
	16'h1280 : data <= 32'h13020000;
	16'h1281 : data <= 32'h93001000;
	16'h1282 : data <= 32'h13017000;
	16'h1283 : data <= 32'hb3912000;
	16'h1284 : data <= 32'h13021200;
	16'h1285 : data <= 32'h93022000;
	16'h1286 : data <= 32'he31652fe;
	16'h1287 : data <= 32'h930e0008;
	16'h1288 : data <= 32'h130ef01b;
	16'h1289 : data <= 32'h6384d101;
	16'h128a : data <= 32'h6f30c002;
	16'h128b : data <= 32'h13020000;
	16'h128c : data <= 32'h93001000;
	16'h128d : data <= 32'h1301e000;
	16'h128e : data <= 32'h13000000;
	16'h128f : data <= 32'hb3912000;
	16'h1290 : data <= 32'h13021200;
	16'h1291 : data <= 32'h93022000;
	16'h1292 : data <= 32'he31452fe;
	16'h1293 : data <= 32'hb74e0000;
	16'h1294 : data <= 32'h130e001c;
	16'h1295 : data <= 32'h6384d101;
	16'h1296 : data <= 32'h6f20d07f;
	16'h1297 : data <= 32'h13020000;
	16'h1298 : data <= 32'h93001000;
	16'h1299 : data <= 32'h1301f001;
	16'h129a : data <= 32'h13000000;
	16'h129b : data <= 32'h13000000;
	16'h129c : data <= 32'hb3912000;
	16'h129d : data <= 32'h13021200;
	16'h129e : data <= 32'h93022000;
	16'h129f : data <= 32'he31252fe;
	16'h12a0 : data <= 32'hb70e0080;
	16'h12a1 : data <= 32'h130e101c;
	16'h12a2 : data <= 32'h6384d101;
	16'h12a3 : data <= 32'h6f20907c;
	16'h12a4 : data <= 32'h13020000;
	16'h12a5 : data <= 32'h93001000;
	16'h12a6 : data <= 32'h13000000;
	16'h12a7 : data <= 32'h13017000;
	16'h12a8 : data <= 32'hb3912000;
	16'h12a9 : data <= 32'h13021200;
	16'h12aa : data <= 32'h93022000;
	16'h12ab : data <= 32'he31452fe;
	16'h12ac : data <= 32'h930e0008;
	16'h12ad : data <= 32'h130e201c;
	16'h12ae : data <= 32'h6384d101;
	16'h12af : data <= 32'h6f209079;
	16'h12b0 : data <= 32'h13020000;
	16'h12b1 : data <= 32'h93001000;
	16'h12b2 : data <= 32'h13000000;
	16'h12b3 : data <= 32'h1301e000;
	16'h12b4 : data <= 32'h13000000;
	16'h12b5 : data <= 32'hb3912000;
	16'h12b6 : data <= 32'h13021200;
	16'h12b7 : data <= 32'h93022000;
	16'h12b8 : data <= 32'he31252fe;
	16'h12b9 : data <= 32'hb74e0000;
	16'h12ba : data <= 32'h130e301c;
	16'h12bb : data <= 32'h6384d101;
	16'h12bc : data <= 32'h6f205076;
	16'h12bd : data <= 32'h13020000;
	16'h12be : data <= 32'h93001000;
	16'h12bf : data <= 32'h13000000;
	16'h12c0 : data <= 32'h13000000;
	16'h12c1 : data <= 32'h1301f001;
	16'h12c2 : data <= 32'hb3912000;
	16'h12c3 : data <= 32'h13021200;
	16'h12c4 : data <= 32'h93022000;
	16'h12c5 : data <= 32'he31252fe;
	16'h12c6 : data <= 32'hb70e0080;
	16'h12c7 : data <= 32'h130e401c;
	16'h12c8 : data <= 32'h6384d101;
	16'h12c9 : data <= 32'h6f201073;
	16'h12ca : data <= 32'h13020000;
	16'h12cb : data <= 32'h13017000;
	16'h12cc : data <= 32'h93001000;
	16'h12cd : data <= 32'hb3912000;
	16'h12ce : data <= 32'h13021200;
	16'h12cf : data <= 32'h93022000;
	16'h12d0 : data <= 32'he31652fe;
	16'h12d1 : data <= 32'h930e0008;
	16'h12d2 : data <= 32'h130e501c;
	16'h12d3 : data <= 32'h6384d101;
	16'h12d4 : data <= 32'h6f205070;
	16'h12d5 : data <= 32'h13020000;
	16'h12d6 : data <= 32'h1301e000;
	16'h12d7 : data <= 32'h93001000;
	16'h12d8 : data <= 32'h13000000;
	16'h12d9 : data <= 32'hb3912000;
	16'h12da : data <= 32'h13021200;
	16'h12db : data <= 32'h93022000;
	16'h12dc : data <= 32'he31452fe;
	16'h12dd : data <= 32'hb74e0000;
	16'h12de : data <= 32'h130e601c;
	16'h12df : data <= 32'h6384d101;
	16'h12e0 : data <= 32'h6f20506d;
	16'h12e1 : data <= 32'h13020000;
	16'h12e2 : data <= 32'h1301f001;
	16'h12e3 : data <= 32'h93001000;
	16'h12e4 : data <= 32'h13000000;
	16'h12e5 : data <= 32'h13000000;
	16'h12e6 : data <= 32'hb3912000;
	16'h12e7 : data <= 32'h13021200;
	16'h12e8 : data <= 32'h93022000;
	16'h12e9 : data <= 32'he31252fe;
	16'h12ea : data <= 32'hb70e0080;
	16'h12eb : data <= 32'h130e701c;
	16'h12ec : data <= 32'h6384d101;
	16'h12ed : data <= 32'h6f20106a;
	16'h12ee : data <= 32'h13020000;
	16'h12ef : data <= 32'h13017000;
	16'h12f0 : data <= 32'h13000000;
	16'h12f1 : data <= 32'h93001000;
	16'h12f2 : data <= 32'hb3912000;
	16'h12f3 : data <= 32'h13021200;
	16'h12f4 : data <= 32'h93022000;
	16'h12f5 : data <= 32'he31452fe;
	16'h12f6 : data <= 32'h930e0008;
	16'h12f7 : data <= 32'h130e801c;
	16'h12f8 : data <= 32'h6384d101;
	16'h12f9 : data <= 32'h6f201067;
	16'h12fa : data <= 32'h13020000;
	16'h12fb : data <= 32'h1301e000;
	16'h12fc : data <= 32'h13000000;
	16'h12fd : data <= 32'h93001000;
	16'h12fe : data <= 32'h13000000;
	16'h12ff : data <= 32'hb3912000;
	16'h1300 : data <= 32'h13021200;
	16'h1301 : data <= 32'h93022000;
	16'h1302 : data <= 32'he31252fe;
	16'h1303 : data <= 32'hb74e0000;
	16'h1304 : data <= 32'h130e901c;
	16'h1305 : data <= 32'h6384d101;
	16'h1306 : data <= 32'h6f20d063;
	16'h1307 : data <= 32'h13020000;
	16'h1308 : data <= 32'h1301f001;
	16'h1309 : data <= 32'h13000000;
	16'h130a : data <= 32'h13000000;
	16'h130b : data <= 32'h93001000;
	16'h130c : data <= 32'hb3912000;
	16'h130d : data <= 32'h13021200;
	16'h130e : data <= 32'h93022000;
	16'h130f : data <= 32'he31252fe;
	16'h1310 : data <= 32'hb70e0080;
	16'h1311 : data <= 32'h130ea01c;
	16'h1312 : data <= 32'h6384d101;
	16'h1313 : data <= 32'h6f209060;
	16'h1314 : data <= 32'h9300f000;
	16'h1315 : data <= 32'h33111000;
	16'h1316 : data <= 32'h930e0000;
	16'h1317 : data <= 32'h130eb01c;
	16'h1318 : data <= 32'h6304d101;
	16'h1319 : data <= 32'h6f20105f;
	16'h131a : data <= 32'h93000002;
	16'h131b : data <= 32'h33910000;
	16'h131c : data <= 32'h930e0002;
	16'h131d : data <= 32'h130ec01c;
	16'h131e : data <= 32'h6304d101;
	16'h131f : data <= 32'h6f20905d;
	16'h1320 : data <= 32'hb3100000;
	16'h1321 : data <= 32'h930e0000;
	16'h1322 : data <= 32'h130ed01c;
	16'h1323 : data <= 32'h6384d001;
	16'h1324 : data <= 32'h6f20505c;
	16'h1325 : data <= 32'h93000040;
	16'h1326 : data <= 32'h37110000;
	16'h1327 : data <= 32'h13010180;
	16'h1328 : data <= 32'h33902000;
	16'h1329 : data <= 32'h930e0000;
	16'h132a : data <= 32'h130ee01c;
	16'h132b : data <= 32'h6304d001;
	16'h132c : data <= 32'h6f20505a;
	16'h132d : data <= 32'h93001000;
	16'h132e : data <= 32'h93910000;
	16'h132f : data <= 32'h930e1000;
	16'h1330 : data <= 32'h130ef01c;
	16'h1331 : data <= 32'h6384d101;
	16'h1332 : data <= 32'h6f20d058;
	16'h1333 : data <= 32'h93001000;
	16'h1334 : data <= 32'h93911000;
	16'h1335 : data <= 32'h930e2000;
	16'h1336 : data <= 32'h130e001d;
	16'h1337 : data <= 32'h6384d101;
	16'h1338 : data <= 32'h6f205057;
	16'h1339 : data <= 32'h93001000;
	16'h133a : data <= 32'h93917000;
	16'h133b : data <= 32'h930e0008;
	16'h133c : data <= 32'h130e101d;
	16'h133d : data <= 32'h6384d101;
	16'h133e : data <= 32'h6f20d055;
	16'h133f : data <= 32'h93001000;
	16'h1340 : data <= 32'h9391e000;
	16'h1341 : data <= 32'hb74e0000;
	16'h1342 : data <= 32'h130e201d;
	16'h1343 : data <= 32'h6384d101;
	16'h1344 : data <= 32'h6f205054;
	16'h1345 : data <= 32'h93001000;
	16'h1346 : data <= 32'h9391f001;
	16'h1347 : data <= 32'hb70e0080;
	16'h1348 : data <= 32'h130e301d;
	16'h1349 : data <= 32'h6384d101;
	16'h134a : data <= 32'h6f20d052;
	16'h134b : data <= 32'h9300f0ff;
	16'h134c : data <= 32'h93910000;
	16'h134d : data <= 32'h930ef0ff;
	16'h134e : data <= 32'h130e401d;
	16'h134f : data <= 32'h6384d101;
	16'h1350 : data <= 32'h6f205051;
	16'h1351 : data <= 32'h9300f0ff;
	16'h1352 : data <= 32'h93911000;
	16'h1353 : data <= 32'h930ee0ff;
	16'h1354 : data <= 32'h130e501d;
	16'h1355 : data <= 32'h6384d101;
	16'h1356 : data <= 32'h6f20d04f;
	16'h1357 : data <= 32'h9300f0ff;
	16'h1358 : data <= 32'h93917000;
	16'h1359 : data <= 32'h930e00f8;
	16'h135a : data <= 32'h130e601d;
	16'h135b : data <= 32'h6384d101;
	16'h135c : data <= 32'h6f20504e;
	16'h135d : data <= 32'h9300f0ff;
	16'h135e : data <= 32'h9391e000;
	16'h135f : data <= 32'hb7ceffff;
	16'h1360 : data <= 32'h130e701d;
	16'h1361 : data <= 32'h6384d101;
	16'h1362 : data <= 32'h6f20d04c;
	16'h1363 : data <= 32'h9300f0ff;
	16'h1364 : data <= 32'h9391f001;
	16'h1365 : data <= 32'hb70e0080;
	16'h1366 : data <= 32'h130e801d;
	16'h1367 : data <= 32'h6384d101;
	16'h1368 : data <= 32'h6f20504b;
	16'h1369 : data <= 32'hb7202121;
	16'h136a : data <= 32'h93801012;
	16'h136b : data <= 32'h93910000;
	16'h136c : data <= 32'hb72e2121;
	16'h136d : data <= 32'h938e1e12;
	16'h136e : data <= 32'h130e901d;
	16'h136f : data <= 32'h6384d101;
	16'h1370 : data <= 32'h6f205049;
	16'h1371 : data <= 32'hb7202121;
	16'h1372 : data <= 32'h93801012;
	16'h1373 : data <= 32'h93911000;
	16'h1374 : data <= 32'hb74e4242;
	16'h1375 : data <= 32'h938e2e24;
	16'h1376 : data <= 32'h130ea01d;
	16'h1377 : data <= 32'h6384d101;
	16'h1378 : data <= 32'h6f205047;
	16'h1379 : data <= 32'hb7202121;
	16'h137a : data <= 32'h93801012;
	16'h137b : data <= 32'h93917000;
	16'h137c : data <= 32'hb79e9090;
	16'h137d : data <= 32'h938e0e08;
	16'h137e : data <= 32'h130eb01d;
	16'h137f : data <= 32'h6384d101;
	16'h1380 : data <= 32'h6f205045;
	16'h1381 : data <= 32'hb7202121;
	16'h1382 : data <= 32'h93801012;
	16'h1383 : data <= 32'h9391e000;
	16'h1384 : data <= 32'hb74e4848;
	16'h1385 : data <= 32'h130ec01d;
	16'h1386 : data <= 32'h6384d101;
	16'h1387 : data <= 32'h6f209043;
	16'h1388 : data <= 32'hb7202121;
	16'h1389 : data <= 32'h93801012;
	16'h138a : data <= 32'h9391f001;
	16'h138b : data <= 32'hb70e0080;
	16'h138c : data <= 32'h130ed01d;
	16'h138d : data <= 32'h6384d101;
	16'h138e : data <= 32'h6f20d041;
	16'h138f : data <= 32'h93001000;
	16'h1390 : data <= 32'h93907000;
	16'h1391 : data <= 32'h930e0008;
	16'h1392 : data <= 32'h130ee01d;
	16'h1393 : data <= 32'h6384d001;
	16'h1394 : data <= 32'h6f205040;
	16'h1395 : data <= 32'h13020000;
	16'h1396 : data <= 32'h93001000;
	16'h1397 : data <= 32'h93917000;
	16'h1398 : data <= 32'h13830100;
	16'h1399 : data <= 32'h13021200;
	16'h139a : data <= 32'h93022000;
	16'h139b : data <= 32'he31652fe;
	16'h139c : data <= 32'h930e0008;
	16'h139d : data <= 32'h130ef01d;
	16'h139e : data <= 32'h6304d301;
	16'h139f : data <= 32'h6f20903d;
	16'h13a0 : data <= 32'h13020000;
	16'h13a1 : data <= 32'h93001000;
	16'h13a2 : data <= 32'h9391e000;
	16'h13a3 : data <= 32'h13000000;
	16'h13a4 : data <= 32'h13830100;
	16'h13a5 : data <= 32'h13021200;
	16'h13a6 : data <= 32'h93022000;
	16'h13a7 : data <= 32'he31452fe;
	16'h13a8 : data <= 32'hb74e0000;
	16'h13a9 : data <= 32'h130e001e;
	16'h13aa : data <= 32'h6304d301;
	16'h13ab : data <= 32'h6f20903a;
	16'h13ac : data <= 32'h13020000;
	16'h13ad : data <= 32'h93001000;
	16'h13ae : data <= 32'h9391f001;
	16'h13af : data <= 32'h13000000;
	16'h13b0 : data <= 32'h13000000;
	16'h13b1 : data <= 32'h13830100;
	16'h13b2 : data <= 32'h13021200;
	16'h13b3 : data <= 32'h93022000;
	16'h13b4 : data <= 32'he31252fe;
	16'h13b5 : data <= 32'hb70e0080;
	16'h13b6 : data <= 32'h130e101e;
	16'h13b7 : data <= 32'h6304d301;
	16'h13b8 : data <= 32'h6f205037;
	16'h13b9 : data <= 32'h13020000;
	16'h13ba : data <= 32'h93001000;
	16'h13bb : data <= 32'h93917000;
	16'h13bc : data <= 32'h13021200;
	16'h13bd : data <= 32'h93022000;
	16'h13be : data <= 32'he31852fe;
	16'h13bf : data <= 32'h930e0008;
	16'h13c0 : data <= 32'h130e201e;
	16'h13c1 : data <= 32'h6384d101;
	16'h13c2 : data <= 32'h6f20d034;
	16'h13c3 : data <= 32'h13020000;
	16'h13c4 : data <= 32'h93001000;
	16'h13c5 : data <= 32'h13000000;
	16'h13c6 : data <= 32'h9391e000;
	16'h13c7 : data <= 32'h13021200;
	16'h13c8 : data <= 32'h93022000;
	16'h13c9 : data <= 32'he31652fe;
	16'h13ca : data <= 32'hb74e0000;
	16'h13cb : data <= 32'h130e301e;
	16'h13cc : data <= 32'h6384d101;
	16'h13cd : data <= 32'h6f201032;
	16'h13ce : data <= 32'h13020000;
	16'h13cf : data <= 32'h93001000;
	16'h13d0 : data <= 32'h13000000;
	16'h13d1 : data <= 32'h13000000;
	16'h13d2 : data <= 32'h9391f001;
	16'h13d3 : data <= 32'h13021200;
	16'h13d4 : data <= 32'h93022000;
	16'h13d5 : data <= 32'he31452fe;
	16'h13d6 : data <= 32'hb70e0080;
	16'h13d7 : data <= 32'h130e401e;
	16'h13d8 : data <= 32'h6384d101;
	16'h13d9 : data <= 32'h6f20102f;
	16'h13da : data <= 32'h9310f001;
	16'h13db : data <= 32'h930e0000;
	16'h13dc : data <= 32'h130e501e;
	16'h13dd : data <= 32'h6384d001;
	16'h13de : data <= 32'h6f20d02d;
	16'h13df : data <= 32'h93001002;
	16'h13e0 : data <= 32'h13904001;
	16'h13e1 : data <= 32'h930e0000;
	16'h13e2 : data <= 32'h130e601e;
	16'h13e3 : data <= 32'h6304d001;
	16'h13e4 : data <= 32'h6f20502c;
	16'h13e5 : data <= 32'h93000000;
	16'h13e6 : data <= 32'h13010000;
	16'h13e7 : data <= 32'hb3a12000;
	16'h13e8 : data <= 32'h930e0000;
	16'h13e9 : data <= 32'h130e701e;
	16'h13ea : data <= 32'h6384d101;
	16'h13eb : data <= 32'h6f20902a;
	16'h13ec : data <= 32'h93001000;
	16'h13ed : data <= 32'h13011000;
	16'h13ee : data <= 32'hb3a12000;
	16'h13ef : data <= 32'h930e0000;
	16'h13f0 : data <= 32'h130e801e;
	16'h13f1 : data <= 32'h6384d101;
	16'h13f2 : data <= 32'h6f20d028;
	16'h13f3 : data <= 32'h93003000;
	16'h13f4 : data <= 32'h13017000;
	16'h13f5 : data <= 32'hb3a12000;
	16'h13f6 : data <= 32'h930e1000;
	16'h13f7 : data <= 32'h130e901e;
	16'h13f8 : data <= 32'h6384d101;
	16'h13f9 : data <= 32'h6f201027;
	16'h13fa : data <= 32'h93007000;
	16'h13fb : data <= 32'h13013000;
	16'h13fc : data <= 32'hb3a12000;
	16'h13fd : data <= 32'h930e0000;
	16'h13fe : data <= 32'h130ea01e;
	16'h13ff : data <= 32'h6384d101;
	16'h1400 : data <= 32'h6f205025;
	16'h1401 : data <= 32'h93000000;
	16'h1402 : data <= 32'h3781ffff;
	16'h1403 : data <= 32'hb3a12000;
	16'h1404 : data <= 32'h930e0000;
	16'h1405 : data <= 32'h130eb01e;
	16'h1406 : data <= 32'h6384d101;
	16'h1407 : data <= 32'h6f209023;
	16'h1408 : data <= 32'hb7000080;
	16'h1409 : data <= 32'h13010000;
	16'h140a : data <= 32'hb3a12000;
	16'h140b : data <= 32'h930e1000;
	16'h140c : data <= 32'h130ec01e;
	16'h140d : data <= 32'h6384d101;
	16'h140e : data <= 32'h6f20d021;
	16'h140f : data <= 32'hb7000080;
	16'h1410 : data <= 32'h3781ffff;
	16'h1411 : data <= 32'hb3a12000;
	16'h1412 : data <= 32'h930e1000;
	16'h1413 : data <= 32'h130ed01e;
	16'h1414 : data <= 32'h6384d101;
	16'h1415 : data <= 32'h6f201020;
	16'h1416 : data <= 32'h93000000;
	16'h1417 : data <= 32'h37810000;
	16'h1418 : data <= 32'h1301f1ff;
	16'h1419 : data <= 32'hb3a12000;
	16'h141a : data <= 32'h930e1000;
	16'h141b : data <= 32'h130ee01e;
	16'h141c : data <= 32'h6384d101;
	16'h141d : data <= 32'h6f20101e;
	16'h141e : data <= 32'hb7000080;
	16'h141f : data <= 32'h9380f0ff;
	16'h1420 : data <= 32'h13010000;
	16'h1421 : data <= 32'hb3a12000;
	16'h1422 : data <= 32'h930e0000;
	16'h1423 : data <= 32'h130ef01e;
	16'h1424 : data <= 32'h6384d101;
	16'h1425 : data <= 32'h6f20101c;
	16'h1426 : data <= 32'hb7000080;
	16'h1427 : data <= 32'h9380f0ff;
	16'h1428 : data <= 32'h37810000;
	16'h1429 : data <= 32'h1301f1ff;
	16'h142a : data <= 32'hb3a12000;
	16'h142b : data <= 32'h930e0000;
	16'h142c : data <= 32'h130e001f;
	16'h142d : data <= 32'h6384d101;
	16'h142e : data <= 32'h6f20d019;
	16'h142f : data <= 32'hb7000080;
	16'h1430 : data <= 32'h37810000;
	16'h1431 : data <= 32'h1301f1ff;
	16'h1432 : data <= 32'hb3a12000;
	16'h1433 : data <= 32'h930e1000;
	16'h1434 : data <= 32'h130e101f;
	16'h1435 : data <= 32'h6384d101;
	16'h1436 : data <= 32'h6f20d017;
	16'h1437 : data <= 32'hb7000080;
	16'h1438 : data <= 32'h9380f0ff;
	16'h1439 : data <= 32'h3781ffff;
	16'h143a : data <= 32'hb3a12000;
	16'h143b : data <= 32'h930e0000;
	16'h143c : data <= 32'h130e201f;
	16'h143d : data <= 32'h6384d101;
	16'h143e : data <= 32'h6f20d015;
	16'h143f : data <= 32'h93000000;
	16'h1440 : data <= 32'h1301f0ff;
	16'h1441 : data <= 32'hb3a12000;
	16'h1442 : data <= 32'h930e0000;
	16'h1443 : data <= 32'h130e301f;
	16'h1444 : data <= 32'h6384d101;
	16'h1445 : data <= 32'h6f201014;
	16'h1446 : data <= 32'h9300f0ff;
	16'h1447 : data <= 32'h13011000;
	16'h1448 : data <= 32'hb3a12000;
	16'h1449 : data <= 32'h930e1000;
	16'h144a : data <= 32'h130e401f;
	16'h144b : data <= 32'h6384d101;
	16'h144c : data <= 32'h6f205012;
	16'h144d : data <= 32'h9300f0ff;
	16'h144e : data <= 32'h1301f0ff;
	16'h144f : data <= 32'hb3a12000;
	16'h1450 : data <= 32'h930e0000;
	16'h1451 : data <= 32'h130e501f;
	16'h1452 : data <= 32'h6384d101;
	16'h1453 : data <= 32'h6f209010;
	16'h1454 : data <= 32'h9300e000;
	16'h1455 : data <= 32'h1301d000;
	16'h1456 : data <= 32'hb3a02000;
	16'h1457 : data <= 32'h930e0000;
	16'h1458 : data <= 32'h130e601f;
	16'h1459 : data <= 32'h6384d001;
	16'h145a : data <= 32'h6f20d00e;
	16'h145b : data <= 32'h9300b000;
	16'h145c : data <= 32'h1301d000;
	16'h145d : data <= 32'h33a12000;
	16'h145e : data <= 32'h930e1000;
	16'h145f : data <= 32'h130e701f;
	16'h1460 : data <= 32'h6304d101;
	16'h1461 : data <= 32'h6f20100d;
	16'h1462 : data <= 32'h9300d000;
	16'h1463 : data <= 32'hb3a01000;
	16'h1464 : data <= 32'h930e0000;
	16'h1465 : data <= 32'h130e801f;
	16'h1466 : data <= 32'h6384d001;
	16'h1467 : data <= 32'h6f20900b;
	16'h1468 : data <= 32'h13020000;
	16'h1469 : data <= 32'h9300b000;
	16'h146a : data <= 32'h1301d000;
	16'h146b : data <= 32'hb3a12000;
	16'h146c : data <= 32'h13830100;
	16'h146d : data <= 32'h13021200;
	16'h146e : data <= 32'h93022000;
	16'h146f : data <= 32'he31452fe;
	16'h1470 : data <= 32'h930e1000;
	16'h1471 : data <= 32'h130e901f;
	16'h1472 : data <= 32'h6304d301;
	16'h1473 : data <= 32'h6f209008;
	16'h1474 : data <= 32'h13020000;
	16'h1475 : data <= 32'h9300e000;
	16'h1476 : data <= 32'h1301d000;
	16'h1477 : data <= 32'hb3a12000;
	16'h1478 : data <= 32'h13000000;
	16'h1479 : data <= 32'h13830100;
	16'h147a : data <= 32'h13021200;
	16'h147b : data <= 32'h93022000;
	16'h147c : data <= 32'he31252fe;
	16'h147d : data <= 32'h930e0000;
	16'h147e : data <= 32'h130ea01f;
	16'h147f : data <= 32'h6304d301;
	16'h1480 : data <= 32'h6f205005;
	16'h1481 : data <= 32'h13020000;
	16'h1482 : data <= 32'h9300c000;
	16'h1483 : data <= 32'h1301d000;
	16'h1484 : data <= 32'hb3a12000;
	16'h1485 : data <= 32'h13000000;
	16'h1486 : data <= 32'h13000000;
	16'h1487 : data <= 32'h13830100;
	16'h1488 : data <= 32'h13021200;
	16'h1489 : data <= 32'h93022000;
	16'h148a : data <= 32'he31052fe;
	16'h148b : data <= 32'h930e1000;
	16'h148c : data <= 32'h130eb01f;
	16'h148d : data <= 32'h6304d301;
	16'h148e : data <= 32'h6f20d001;
	16'h148f : data <= 32'h13020000;
	16'h1490 : data <= 32'h9300e000;
	16'h1491 : data <= 32'h1301d000;
	16'h1492 : data <= 32'hb3a12000;
	16'h1493 : data <= 32'h13021200;
	16'h1494 : data <= 32'h93022000;
	16'h1495 : data <= 32'he31652fe;
	16'h1496 : data <= 32'h930e0000;
	16'h1497 : data <= 32'h130ec01f;
	16'h1498 : data <= 32'h6384d101;
	16'h1499 : data <= 32'h6f20007f;
	16'h149a : data <= 32'h13020000;
	16'h149b : data <= 32'h9300b000;
	16'h149c : data <= 32'h1301d000;
	16'h149d : data <= 32'h13000000;
	16'h149e : data <= 32'hb3a12000;
	16'h149f : data <= 32'h13021200;
	16'h14a0 : data <= 32'h93022000;
	16'h14a1 : data <= 32'he31452fe;
	16'h14a2 : data <= 32'h930e1000;
	16'h14a3 : data <= 32'h130ed01f;
	16'h14a4 : data <= 32'h6384d101;
	16'h14a5 : data <= 32'h6f20007c;
	16'h14a6 : data <= 32'h13020000;
	16'h14a7 : data <= 32'h9300f000;
	16'h14a8 : data <= 32'h1301d000;
	16'h14a9 : data <= 32'h13000000;
	16'h14aa : data <= 32'h13000000;
	16'h14ab : data <= 32'hb3a12000;
	16'h14ac : data <= 32'h13021200;
	16'h14ad : data <= 32'h93022000;
	16'h14ae : data <= 32'he31252fe;
	16'h14af : data <= 32'h930e0000;
	16'h14b0 : data <= 32'h130ee01f;
	16'h14b1 : data <= 32'h6384d101;
	16'h14b2 : data <= 32'h6f20c078;
	16'h14b3 : data <= 32'h13020000;
	16'h14b4 : data <= 32'h9300a000;
	16'h14b5 : data <= 32'h13000000;
	16'h14b6 : data <= 32'h1301d000;
	16'h14b7 : data <= 32'hb3a12000;
	16'h14b8 : data <= 32'h13021200;
	16'h14b9 : data <= 32'h93022000;
	16'h14ba : data <= 32'he31452fe;
	16'h14bb : data <= 32'h930e1000;
	16'h14bc : data <= 32'h130ef01f;
	16'h14bd : data <= 32'h6384d101;
	16'h14be : data <= 32'h6f20c075;
	16'h14bf : data <= 32'h13020000;
	16'h14c0 : data <= 32'h93000001;
	16'h14c1 : data <= 32'h13000000;
	16'h14c2 : data <= 32'h1301d000;
	16'h14c3 : data <= 32'h13000000;
	16'h14c4 : data <= 32'hb3a12000;
	16'h14c5 : data <= 32'h13021200;
	16'h14c6 : data <= 32'h93022000;
	16'h14c7 : data <= 32'he31252fe;
	16'h14c8 : data <= 32'h930e0000;
	16'h14c9 : data <= 32'h130e0020;
	16'h14ca : data <= 32'h6384d101;
	16'h14cb : data <= 32'h6f208072;
	16'h14cc : data <= 32'h13020000;
	16'h14cd : data <= 32'h93009000;
	16'h14ce : data <= 32'h13000000;
	16'h14cf : data <= 32'h13000000;
	16'h14d0 : data <= 32'h1301d000;
	16'h14d1 : data <= 32'hb3a12000;
	16'h14d2 : data <= 32'h13021200;
	16'h14d3 : data <= 32'h93022000;
	16'h14d4 : data <= 32'he31252fe;
	16'h14d5 : data <= 32'h930e1000;
	16'h14d6 : data <= 32'h130e1020;
	16'h14d7 : data <= 32'h6384d101;
	16'h14d8 : data <= 32'h6f20406f;
	16'h14d9 : data <= 32'h13020000;
	16'h14da : data <= 32'h1301d000;
	16'h14db : data <= 32'h93001001;
	16'h14dc : data <= 32'hb3a12000;
	16'h14dd : data <= 32'h13021200;
	16'h14de : data <= 32'h93022000;
	16'h14df : data <= 32'he31652fe;
	16'h14e0 : data <= 32'h930e0000;
	16'h14e1 : data <= 32'h130e2020;
	16'h14e2 : data <= 32'h6384d101;
	16'h14e3 : data <= 32'h6f20806c;
	16'h14e4 : data <= 32'h13020000;
	16'h14e5 : data <= 32'h1301d000;
	16'h14e6 : data <= 32'h93008000;
	16'h14e7 : data <= 32'h13000000;
	16'h14e8 : data <= 32'hb3a12000;
	16'h14e9 : data <= 32'h13021200;
	16'h14ea : data <= 32'h93022000;
	16'h14eb : data <= 32'he31452fe;
	16'h14ec : data <= 32'h930e1000;
	16'h14ed : data <= 32'h130e3020;
	16'h14ee : data <= 32'h6384d101;
	16'h14ef : data <= 32'h6f208069;
	16'h14f0 : data <= 32'h13020000;
	16'h14f1 : data <= 32'h1301d000;
	16'h14f2 : data <= 32'h93002001;
	16'h14f3 : data <= 32'h13000000;
	16'h14f4 : data <= 32'h13000000;
	16'h14f5 : data <= 32'hb3a12000;
	16'h14f6 : data <= 32'h13021200;
	16'h14f7 : data <= 32'h93022000;
	16'h14f8 : data <= 32'he31252fe;
	16'h14f9 : data <= 32'h930e0000;
	16'h14fa : data <= 32'h130e4020;
	16'h14fb : data <= 32'h6384d101;
	16'h14fc : data <= 32'h6f204066;
	16'h14fd : data <= 32'h13020000;
	16'h14fe : data <= 32'h1301d000;
	16'h14ff : data <= 32'h13000000;
	16'h1500 : data <= 32'h93007000;
	16'h1501 : data <= 32'hb3a12000;
	16'h1502 : data <= 32'h13021200;
	16'h1503 : data <= 32'h93022000;
	16'h1504 : data <= 32'he31452fe;
	16'h1505 : data <= 32'h930e1000;
	16'h1506 : data <= 32'h130e5020;
	16'h1507 : data <= 32'h6384d101;
	16'h1508 : data <= 32'h6f204063;
	16'h1509 : data <= 32'h13020000;
	16'h150a : data <= 32'h1301d000;
	16'h150b : data <= 32'h13000000;
	16'h150c : data <= 32'h93003001;
	16'h150d : data <= 32'h13000000;
	16'h150e : data <= 32'hb3a12000;
	16'h150f : data <= 32'h13021200;
	16'h1510 : data <= 32'h93022000;
	16'h1511 : data <= 32'he31252fe;
	16'h1512 : data <= 32'h930e0000;
	16'h1513 : data <= 32'h130e6020;
	16'h1514 : data <= 32'h6384d101;
	16'h1515 : data <= 32'h6f200060;
	16'h1516 : data <= 32'h13020000;
	16'h1517 : data <= 32'h1301d000;
	16'h1518 : data <= 32'h13000000;
	16'h1519 : data <= 32'h13000000;
	16'h151a : data <= 32'h93006000;
	16'h151b : data <= 32'hb3a12000;
	16'h151c : data <= 32'h13021200;
	16'h151d : data <= 32'h93022000;
	16'h151e : data <= 32'he31252fe;
	16'h151f : data <= 32'h930e1000;
	16'h1520 : data <= 32'h130e7020;
	16'h1521 : data <= 32'h6384d101;
	16'h1522 : data <= 32'h6f20c05c;
	16'h1523 : data <= 32'h9300f0ff;
	16'h1524 : data <= 32'h33211000;
	16'h1525 : data <= 32'h930e0000;
	16'h1526 : data <= 32'h130e8020;
	16'h1527 : data <= 32'h6304d101;
	16'h1528 : data <= 32'h6f20405b;
	16'h1529 : data <= 32'h9300f0ff;
	16'h152a : data <= 32'h33a10000;
	16'h152b : data <= 32'h930e1000;
	16'h152c : data <= 32'h130e9020;
	16'h152d : data <= 32'h6304d101;
	16'h152e : data <= 32'h6f20c059;
	16'h152f : data <= 32'hb3200000;
	16'h1530 : data <= 32'h930e0000;
	16'h1531 : data <= 32'h130ea020;
	16'h1532 : data <= 32'h6384d001;
	16'h1533 : data <= 32'h6f208058;
	16'h1534 : data <= 32'h93000001;
	16'h1535 : data <= 32'h1301e001;
	16'h1536 : data <= 32'h33a02000;
	16'h1537 : data <= 32'h930e0000;
	16'h1538 : data <= 32'h130eb020;
	16'h1539 : data <= 32'h6304d001;
	16'h153a : data <= 32'h6f20c056;
	16'h153b : data <= 32'h93000000;
	16'h153c : data <= 32'h93a10000;
	16'h153d : data <= 32'h930e0000;
	16'h153e : data <= 32'h130ec020;
	16'h153f : data <= 32'h6384d101;
	16'h1540 : data <= 32'h6f204055;
	16'h1541 : data <= 32'h93001000;
	16'h1542 : data <= 32'h93a11000;
	16'h1543 : data <= 32'h930e0000;
	16'h1544 : data <= 32'h130ed020;
	16'h1545 : data <= 32'h6384d101;
	16'h1546 : data <= 32'h6f20c053;
	16'h1547 : data <= 32'h93003000;
	16'h1548 : data <= 32'h93a17000;
	16'h1549 : data <= 32'h930e1000;
	16'h154a : data <= 32'h130ee020;
	16'h154b : data <= 32'h6384d101;
	16'h154c : data <= 32'h6f204052;
	16'h154d : data <= 32'h93007000;
	16'h154e : data <= 32'h93a13000;
	16'h154f : data <= 32'h930e0000;
	16'h1550 : data <= 32'h130ef020;
	16'h1551 : data <= 32'h6384d101;
	16'h1552 : data <= 32'h6f20c050;
	16'h1553 : data <= 32'h93000000;
	16'h1554 : data <= 32'h93a10080;
	16'h1555 : data <= 32'h930e0000;
	16'h1556 : data <= 32'h130e0021;
	16'h1557 : data <= 32'h6384d101;
	16'h1558 : data <= 32'h6f20404f;
	16'h1559 : data <= 32'hb7000080;
	16'h155a : data <= 32'h93a10000;
	16'h155b : data <= 32'h930e1000;
	16'h155c : data <= 32'h130e1021;
	16'h155d : data <= 32'h6384d101;
	16'h155e : data <= 32'h6f20c04d;
	16'h155f : data <= 32'hb7000080;
	16'h1560 : data <= 32'h93a10080;
	16'h1561 : data <= 32'h930e1000;
	16'h1562 : data <= 32'h130e2021;
	16'h1563 : data <= 32'h6384d101;
	16'h1564 : data <= 32'h6f20404c;
	16'h1565 : data <= 32'h93000000;
	16'h1566 : data <= 32'h93a1f07f;
	16'h1567 : data <= 32'h930e1000;
	16'h1568 : data <= 32'h130e3021;
	16'h1569 : data <= 32'h6384d101;
	16'h156a : data <= 32'h6f20c04a;
	16'h156b : data <= 32'hb7000080;
	16'h156c : data <= 32'h9380f0ff;
	16'h156d : data <= 32'h93a10000;
	16'h156e : data <= 32'h930e0000;
	16'h156f : data <= 32'h130e4021;
	16'h1570 : data <= 32'h6384d101;
	16'h1571 : data <= 32'h6f200049;
	16'h1572 : data <= 32'hb7000080;
	16'h1573 : data <= 32'h9380f0ff;
	16'h1574 : data <= 32'h93a1f07f;
	16'h1575 : data <= 32'h930e0000;
	16'h1576 : data <= 32'h130e5021;
	16'h1577 : data <= 32'h6384d101;
	16'h1578 : data <= 32'h6f204047;
	16'h1579 : data <= 32'hb7000080;
	16'h157a : data <= 32'h93a1f07f;
	16'h157b : data <= 32'h930e1000;
	16'h157c : data <= 32'h130e6021;
	16'h157d : data <= 32'h6384d101;
	16'h157e : data <= 32'h6f20c045;
	16'h157f : data <= 32'hb7000080;
	16'h1580 : data <= 32'h9380f0ff;
	16'h1581 : data <= 32'h93a10080;
	16'h1582 : data <= 32'h930e0000;
	16'h1583 : data <= 32'h130e7021;
	16'h1584 : data <= 32'h6384d101;
	16'h1585 : data <= 32'h6f200044;
	16'h1586 : data <= 32'h93000000;
	16'h1587 : data <= 32'h93a1f0ff;
	16'h1588 : data <= 32'h930e0000;
	16'h1589 : data <= 32'h130e8021;
	16'h158a : data <= 32'h6384d101;
	16'h158b : data <= 32'h6f208042;
	16'h158c : data <= 32'h9300f0ff;
	16'h158d : data <= 32'h93a11000;
	16'h158e : data <= 32'h930e1000;
	16'h158f : data <= 32'h130e9021;
	16'h1590 : data <= 32'h6384d101;
	16'h1591 : data <= 32'h6f200041;
	16'h1592 : data <= 32'h9300f0ff;
	16'h1593 : data <= 32'h93a1f0ff;
	16'h1594 : data <= 32'h930e0000;
	16'h1595 : data <= 32'h130ea021;
	16'h1596 : data <= 32'h6384d101;
	16'h1597 : data <= 32'h6f20803f;
	16'h1598 : data <= 32'h9300b000;
	16'h1599 : data <= 32'h93b0d000;
	16'h159a : data <= 32'h930e1000;
	16'h159b : data <= 32'h130eb021;
	16'h159c : data <= 32'h6384d001;
	16'h159d : data <= 32'h6f20003e;
	16'h159e : data <= 32'h13020000;
	16'h159f : data <= 32'h9300f000;
	16'h15a0 : data <= 32'h93a1a000;
	16'h15a1 : data <= 32'h13830100;
	16'h15a2 : data <= 32'h13021200;
	16'h15a3 : data <= 32'h93022000;
	16'h15a4 : data <= 32'he31652fe;
	16'h15a5 : data <= 32'h930e0000;
	16'h15a6 : data <= 32'h130ec021;
	16'h15a7 : data <= 32'h6304d301;
	16'h15a8 : data <= 32'h6f20403b;
	16'h15a9 : data <= 32'h13020000;
	16'h15aa : data <= 32'h9300a000;
	16'h15ab : data <= 32'h93a10001;
	16'h15ac : data <= 32'h13000000;
	16'h15ad : data <= 32'h13830100;
	16'h15ae : data <= 32'h13021200;
	16'h15af : data <= 32'h93022000;
	16'h15b0 : data <= 32'he31452fe;
	16'h15b1 : data <= 32'h930e1000;
	16'h15b2 : data <= 32'h130ed021;
	16'h15b3 : data <= 32'h6304d301;
	16'h15b4 : data <= 32'h6f204038;
	16'h15b5 : data <= 32'h13020000;
	16'h15b6 : data <= 32'h93000001;
	16'h15b7 : data <= 32'h93a19000;
	16'h15b8 : data <= 32'h13000000;
	16'h15b9 : data <= 32'h13000000;
	16'h15ba : data <= 32'h13830100;
	16'h15bb : data <= 32'h13021200;
	16'h15bc : data <= 32'h93022000;
	16'h15bd : data <= 32'he31252fe;
	16'h15be : data <= 32'h930e0000;
	16'h15bf : data <= 32'h130ee021;
	16'h15c0 : data <= 32'h6304d301;
	16'h15c1 : data <= 32'h6f200035;
	16'h15c2 : data <= 32'h13020000;
	16'h15c3 : data <= 32'h9300b000;
	16'h15c4 : data <= 32'h93a1f000;
	16'h15c5 : data <= 32'h13021200;
	16'h15c6 : data <= 32'h93022000;
	16'h15c7 : data <= 32'he31852fe;
	16'h15c8 : data <= 32'h930e1000;
	16'h15c9 : data <= 32'h130ef021;
	16'h15ca : data <= 32'h6384d101;
	16'h15cb : data <= 32'h6f208032;
	16'h15cc : data <= 32'h13020000;
	16'h15cd : data <= 32'h93001001;
	16'h15ce : data <= 32'h13000000;
	16'h15cf : data <= 32'h93a18000;
	16'h15d0 : data <= 32'h13021200;
	16'h15d1 : data <= 32'h93022000;
	16'h15d2 : data <= 32'he31652fe;
	16'h15d3 : data <= 32'h930e0000;
	16'h15d4 : data <= 32'h130e0022;
	16'h15d5 : data <= 32'h6384d101;
	16'h15d6 : data <= 32'h6f20c02f;
	16'h15d7 : data <= 32'h13020000;
	16'h15d8 : data <= 32'h9300c000;
	16'h15d9 : data <= 32'h13000000;
	16'h15da : data <= 32'h13000000;
	16'h15db : data <= 32'h93a1e000;
	16'h15dc : data <= 32'h13021200;
	16'h15dd : data <= 32'h93022000;
	16'h15de : data <= 32'he31452fe;
	16'h15df : data <= 32'h930e1000;
	16'h15e0 : data <= 32'h130e1022;
	16'h15e1 : data <= 32'h6384d101;
	16'h15e2 : data <= 32'h6f20c02c;
	16'h15e3 : data <= 32'h9320f0ff;
	16'h15e4 : data <= 32'h930e0000;
	16'h15e5 : data <= 32'h130e2022;
	16'h15e6 : data <= 32'h6384d001;
	16'h15e7 : data <= 32'h6f20802b;
	16'h15e8 : data <= 32'hb700ff00;
	16'h15e9 : data <= 32'h9380f00f;
	16'h15ea : data <= 32'h13a0f0ff;
	16'h15eb : data <= 32'h930e0000;
	16'h15ec : data <= 32'h130e3022;
	16'h15ed : data <= 32'h6304d001;
	16'h15ee : data <= 32'h6f20c029;
	16'h15ef : data <= 32'hb7000080;
	16'h15f0 : data <= 32'h13010000;
	16'h15f1 : data <= 32'hb3d12040;
	16'h15f2 : data <= 32'hb70e0080;
	16'h15f3 : data <= 32'h130e4022;
	16'h15f4 : data <= 32'h6384d101;
	16'h15f5 : data <= 32'h6f200028;
	16'h15f6 : data <= 32'hb7000080;
	16'h15f7 : data <= 32'h13011000;
	16'h15f8 : data <= 32'hb3d12040;
	16'h15f9 : data <= 32'hb70e00c0;
	16'h15fa : data <= 32'h130e5022;
	16'h15fb : data <= 32'h6384d101;
	16'h15fc : data <= 32'h6f204026;
	16'h15fd : data <= 32'hb7000080;
	16'h15fe : data <= 32'h13017000;
	16'h15ff : data <= 32'hb3d12040;
	16'h1600 : data <= 32'hb70e00ff;
	16'h1601 : data <= 32'h130e6022;
	16'h1602 : data <= 32'h6384d101;
	16'h1603 : data <= 32'h6f208024;
	16'h1604 : data <= 32'hb7000080;
	16'h1605 : data <= 32'h1301e000;
	16'h1606 : data <= 32'hb3d12040;
	16'h1607 : data <= 32'hb70efeff;
	16'h1608 : data <= 32'h130e7022;
	16'h1609 : data <= 32'h6384d101;
	16'h160a : data <= 32'h6f20c022;
	16'h160b : data <= 32'hb7000080;
	16'h160c : data <= 32'h93801000;
	16'h160d : data <= 32'h1301f001;
	16'h160e : data <= 32'hb3d12040;
	16'h160f : data <= 32'h930ef0ff;
	16'h1610 : data <= 32'h130e8022;
	16'h1611 : data <= 32'h6384d101;
	16'h1612 : data <= 32'h6f20c020;
	16'h1613 : data <= 32'hb7000080;
	16'h1614 : data <= 32'h9380f0ff;
	16'h1615 : data <= 32'h13010000;
	16'h1616 : data <= 32'hb3d12040;
	16'h1617 : data <= 32'hb70e0080;
	16'h1618 : data <= 32'h938efeff;
	16'h1619 : data <= 32'h130e9022;
	16'h161a : data <= 32'h6384d101;
	16'h161b : data <= 32'h6f20801e;
	16'h161c : data <= 32'hb7000080;
	16'h161d : data <= 32'h9380f0ff;
	16'h161e : data <= 32'h13011000;
	16'h161f : data <= 32'hb3d12040;
	16'h1620 : data <= 32'hb70e0040;
	16'h1621 : data <= 32'h938efeff;
	16'h1622 : data <= 32'h130ea022;
	16'h1623 : data <= 32'h6384d101;
	16'h1624 : data <= 32'h6f20401c;
	16'h1625 : data <= 32'hb7000080;
	16'h1626 : data <= 32'h9380f0ff;
	16'h1627 : data <= 32'h13017000;
	16'h1628 : data <= 32'hb3d12040;
	16'h1629 : data <= 32'hb70e0001;
	16'h162a : data <= 32'h938efeff;
	16'h162b : data <= 32'h130eb022;
	16'h162c : data <= 32'h6384d101;
	16'h162d : data <= 32'h6f20001a;
	16'h162e : data <= 32'hb7000080;
	16'h162f : data <= 32'h9380f0ff;
	16'h1630 : data <= 32'h1301e000;
	16'h1631 : data <= 32'hb3d12040;
	16'h1632 : data <= 32'hb70e0200;
	16'h1633 : data <= 32'h938efeff;
	16'h1634 : data <= 32'h130ec022;
	16'h1635 : data <= 32'h6384d101;
	16'h1636 : data <= 32'h6f20c017;
	16'h1637 : data <= 32'hb7000080;
	16'h1638 : data <= 32'h9380f0ff;
	16'h1639 : data <= 32'h1301f001;
	16'h163a : data <= 32'hb3d12040;
	16'h163b : data <= 32'h930e0000;
	16'h163c : data <= 32'h130ed022;
	16'h163d : data <= 32'h6384d101;
	16'h163e : data <= 32'h6f20c015;
	16'h163f : data <= 32'hb7808181;
	16'h1640 : data <= 32'h93801018;
	16'h1641 : data <= 32'h13010000;
	16'h1642 : data <= 32'hb3d12040;
	16'h1643 : data <= 32'hb78e8181;
	16'h1644 : data <= 32'h938e1e18;
	16'h1645 : data <= 32'h130ee022;
	16'h1646 : data <= 32'h6384d101;
	16'h1647 : data <= 32'h6f208013;
	16'h1648 : data <= 32'hb7808181;
	16'h1649 : data <= 32'h93801018;
	16'h164a : data <= 32'h13011000;
	16'h164b : data <= 32'hb3d12040;
	16'h164c : data <= 32'hb7cec0c0;
	16'h164d : data <= 32'h938e0e0c;
	16'h164e : data <= 32'h130ef022;
	16'h164f : data <= 32'h6384d101;
	16'h1650 : data <= 32'h6f204011;
	16'h1651 : data <= 32'hb7808181;
	16'h1652 : data <= 32'h93801018;
	16'h1653 : data <= 32'h13017000;
	16'h1654 : data <= 32'hb3d12040;
	16'h1655 : data <= 32'hb70e03ff;
	16'h1656 : data <= 32'h938e3e30;
	16'h1657 : data <= 32'h130e0023;
	16'h1658 : data <= 32'h6384d101;
	16'h1659 : data <= 32'h6f20000f;
	16'h165a : data <= 32'hb7808181;
	16'h165b : data <= 32'h93801018;
	16'h165c : data <= 32'h1301e000;
	16'h165d : data <= 32'hb3d12040;
	16'h165e : data <= 32'hb70efeff;
	16'h165f : data <= 32'h938e6e60;
	16'h1660 : data <= 32'h130e1023;
	16'h1661 : data <= 32'h6384d101;
	16'h1662 : data <= 32'h6f20c00c;
	16'h1663 : data <= 32'hb7808181;
	16'h1664 : data <= 32'h93801018;
	16'h1665 : data <= 32'h1301f001;
	16'h1666 : data <= 32'hb3d12040;
	16'h1667 : data <= 32'h930ef0ff;
	16'h1668 : data <= 32'h130e2023;
	16'h1669 : data <= 32'h6384d101;
	16'h166a : data <= 32'h6f20c00a;
	16'h166b : data <= 32'hb7808181;
	16'h166c : data <= 32'h93801018;
	16'h166d : data <= 32'h130100fc;
	16'h166e : data <= 32'hb3d12040;
	16'h166f : data <= 32'hb78e8181;
	16'h1670 : data <= 32'h938e1e18;
	16'h1671 : data <= 32'h130e3023;
	16'h1672 : data <= 32'h6384d101;
	16'h1673 : data <= 32'h6f208008;
	16'h1674 : data <= 32'hb7808181;
	16'h1675 : data <= 32'h93801018;
	16'h1676 : data <= 32'h130110fc;
	16'h1677 : data <= 32'hb3d12040;
	16'h1678 : data <= 32'hb7cec0c0;
	16'h1679 : data <= 32'h938e0e0c;
	16'h167a : data <= 32'h130e4023;
	16'h167b : data <= 32'h6384d101;
	16'h167c : data <= 32'h6f204006;
	16'h167d : data <= 32'hb7808181;
	16'h167e : data <= 32'h93801018;
	16'h167f : data <= 32'h130170fc;
	16'h1680 : data <= 32'hb3d12040;
	16'h1681 : data <= 32'hb70e03ff;
	16'h1682 : data <= 32'h938e3e30;
	16'h1683 : data <= 32'h130e5023;
	16'h1684 : data <= 32'h6384d101;
	16'h1685 : data <= 32'h6f200004;
	16'h1686 : data <= 32'hb7808181;
	16'h1687 : data <= 32'h93801018;
	16'h1688 : data <= 32'h1301e0fc;
	16'h1689 : data <= 32'hb3d12040;
	16'h168a : data <= 32'hb70efeff;
	16'h168b : data <= 32'h938e6e60;
	16'h168c : data <= 32'h130e6023;
	16'h168d : data <= 32'h6384d101;
	16'h168e : data <= 32'h6f20c001;
	16'h168f : data <= 32'hb7808181;
	16'h1690 : data <= 32'h93801018;
	16'h1691 : data <= 32'h1301f0ff;
	16'h1692 : data <= 32'hb3d12040;
	16'h1693 : data <= 32'h930ef0ff;
	16'h1694 : data <= 32'h130e7023;
	16'h1695 : data <= 32'h6384d101;
	16'h1696 : data <= 32'h6f10d07f;
	16'h1697 : data <= 32'hb7000080;
	16'h1698 : data <= 32'h13017000;
	16'h1699 : data <= 32'hb3d02040;
	16'h169a : data <= 32'hb70e00ff;
	16'h169b : data <= 32'h130e8023;
	16'h169c : data <= 32'h6384d001;
	16'h169d : data <= 32'h6f10107e;
	16'h169e : data <= 32'hb7000080;
	16'h169f : data <= 32'h1301e000;
	16'h16a0 : data <= 32'h33d12040;
	16'h16a1 : data <= 32'hb70efeff;
	16'h16a2 : data <= 32'h130e9023;
	16'h16a3 : data <= 32'h6304d101;
	16'h16a4 : data <= 32'h6f10507c;
	16'h16a5 : data <= 32'h93007000;
	16'h16a6 : data <= 32'hb3d01040;
	16'h16a7 : data <= 32'h930e0000;
	16'h16a8 : data <= 32'h130ea023;
	16'h16a9 : data <= 32'h6384d001;
	16'h16aa : data <= 32'h6f10d07a;
	16'h16ab : data <= 32'h13020000;
	16'h16ac : data <= 32'hb7000080;
	16'h16ad : data <= 32'h13017000;
	16'h16ae : data <= 32'hb3d12040;
	16'h16af : data <= 32'h13830100;
	16'h16b0 : data <= 32'h13021200;
	16'h16b1 : data <= 32'h93022000;
	16'h16b2 : data <= 32'he31452fe;
	16'h16b3 : data <= 32'hb70e00ff;
	16'h16b4 : data <= 32'h130eb023;
	16'h16b5 : data <= 32'h6304d301;
	16'h16b6 : data <= 32'h6f10d077;
	16'h16b7 : data <= 32'h13020000;
	16'h16b8 : data <= 32'hb7000080;
	16'h16b9 : data <= 32'h1301e000;
	16'h16ba : data <= 32'hb3d12040;
	16'h16bb : data <= 32'h13000000;
	16'h16bc : data <= 32'h13830100;
	16'h16bd : data <= 32'h13021200;
	16'h16be : data <= 32'h93022000;
	16'h16bf : data <= 32'he31252fe;
	16'h16c0 : data <= 32'hb70efeff;
	16'h16c1 : data <= 32'h130ec023;
	16'h16c2 : data <= 32'h6304d301;
	16'h16c3 : data <= 32'h6f109074;
	16'h16c4 : data <= 32'h13020000;
	16'h16c5 : data <= 32'hb7000080;
	16'h16c6 : data <= 32'h1301f001;
	16'h16c7 : data <= 32'hb3d12040;
	16'h16c8 : data <= 32'h13000000;
	16'h16c9 : data <= 32'h13000000;
	16'h16ca : data <= 32'h13830100;
	16'h16cb : data <= 32'h13021200;
	16'h16cc : data <= 32'h93022000;
	16'h16cd : data <= 32'he31052fe;
	16'h16ce : data <= 32'h930ef0ff;
	16'h16cf : data <= 32'h130ed023;
	16'h16d0 : data <= 32'h6304d301;
	16'h16d1 : data <= 32'h6f101071;
	16'h16d2 : data <= 32'h13020000;
	16'h16d3 : data <= 32'hb7000080;
	16'h16d4 : data <= 32'h13017000;
	16'h16d5 : data <= 32'hb3d12040;
	16'h16d6 : data <= 32'h13021200;
	16'h16d7 : data <= 32'h93022000;
	16'h16d8 : data <= 32'he31652fe;
	16'h16d9 : data <= 32'hb70e00ff;
	16'h16da : data <= 32'h130ee023;
	16'h16db : data <= 32'h6384d101;
	16'h16dc : data <= 32'h6f10506e;
	16'h16dd : data <= 32'h13020000;
	16'h16de : data <= 32'hb7000080;
	16'h16df : data <= 32'h1301e000;
	16'h16e0 : data <= 32'h13000000;
	16'h16e1 : data <= 32'hb3d12040;
	16'h16e2 : data <= 32'h13021200;
	16'h16e3 : data <= 32'h93022000;
	16'h16e4 : data <= 32'he31452fe;
	16'h16e5 : data <= 32'hb70efeff;
	16'h16e6 : data <= 32'h130ef023;
	16'h16e7 : data <= 32'h6384d101;
	16'h16e8 : data <= 32'h6f10506b;
	16'h16e9 : data <= 32'h13020000;
	16'h16ea : data <= 32'hb7000080;
	16'h16eb : data <= 32'h1301f001;
	16'h16ec : data <= 32'h13000000;
	16'h16ed : data <= 32'h13000000;
	16'h16ee : data <= 32'hb3d12040;
	16'h16ef : data <= 32'h13021200;
	16'h16f0 : data <= 32'h93022000;
	16'h16f1 : data <= 32'he31252fe;
	16'h16f2 : data <= 32'h930ef0ff;
	16'h16f3 : data <= 32'h130e0024;
	16'h16f4 : data <= 32'h6384d101;
	16'h16f5 : data <= 32'h6f101068;
	16'h16f6 : data <= 32'h13020000;
	16'h16f7 : data <= 32'hb7000080;
	16'h16f8 : data <= 32'h13000000;
	16'h16f9 : data <= 32'h13017000;
	16'h16fa : data <= 32'hb3d12040;
	16'h16fb : data <= 32'h13021200;
	16'h16fc : data <= 32'h93022000;
	16'h16fd : data <= 32'he31452fe;
	16'h16fe : data <= 32'hb70e00ff;
	16'h16ff : data <= 32'h130e1024;
	16'h1700 : data <= 32'h6384d101;
	16'h1701 : data <= 32'h6f101065;
	16'h1702 : data <= 32'h13020000;
	16'h1703 : data <= 32'hb7000080;
	16'h1704 : data <= 32'h13000000;
	16'h1705 : data <= 32'h1301e000;
	16'h1706 : data <= 32'h13000000;
	16'h1707 : data <= 32'hb3d12040;
	16'h1708 : data <= 32'h13021200;
	16'h1709 : data <= 32'h93022000;
	16'h170a : data <= 32'he31252fe;
	16'h170b : data <= 32'hb70efeff;
	16'h170c : data <= 32'h130e2024;
	16'h170d : data <= 32'h6384d101;
	16'h170e : data <= 32'h6f10d061;
	16'h170f : data <= 32'h13020000;
	16'h1710 : data <= 32'hb7000080;
	16'h1711 : data <= 32'h13000000;
	16'h1712 : data <= 32'h13000000;
	16'h1713 : data <= 32'h1301f001;
	16'h1714 : data <= 32'hb3d12040;
	16'h1715 : data <= 32'h13021200;
	16'h1716 : data <= 32'h93022000;
	16'h1717 : data <= 32'he31252fe;
	16'h1718 : data <= 32'h930ef0ff;
	16'h1719 : data <= 32'h130e3024;
	16'h171a : data <= 32'h6384d101;
	16'h171b : data <= 32'h6f10905e;
	16'h171c : data <= 32'h13020000;
	16'h171d : data <= 32'h13017000;
	16'h171e : data <= 32'hb7000080;
	16'h171f : data <= 32'hb3d12040;
	16'h1720 : data <= 32'h13021200;
	16'h1721 : data <= 32'h93022000;
	16'h1722 : data <= 32'he31652fe;
	16'h1723 : data <= 32'hb70e00ff;
	16'h1724 : data <= 32'h130e4024;
	16'h1725 : data <= 32'h6384d101;
	16'h1726 : data <= 32'h6f10d05b;
	16'h1727 : data <= 32'h13020000;
	16'h1728 : data <= 32'h1301e000;
	16'h1729 : data <= 32'hb7000080;
	16'h172a : data <= 32'h13000000;
	16'h172b : data <= 32'hb3d12040;
	16'h172c : data <= 32'h13021200;
	16'h172d : data <= 32'h93022000;
	16'h172e : data <= 32'he31452fe;
	16'h172f : data <= 32'hb70efeff;
	16'h1730 : data <= 32'h130e5024;
	16'h1731 : data <= 32'h6384d101;
	16'h1732 : data <= 32'h6f10d058;
	16'h1733 : data <= 32'h13020000;
	16'h1734 : data <= 32'h1301f001;
	16'h1735 : data <= 32'hb7000080;
	16'h1736 : data <= 32'h13000000;
	16'h1737 : data <= 32'h13000000;
	16'h1738 : data <= 32'hb3d12040;
	16'h1739 : data <= 32'h13021200;
	16'h173a : data <= 32'h93022000;
	16'h173b : data <= 32'he31252fe;
	16'h173c : data <= 32'h930ef0ff;
	16'h173d : data <= 32'h130e6024;
	16'h173e : data <= 32'h6384d101;
	16'h173f : data <= 32'h6f109055;
	16'h1740 : data <= 32'h13020000;
	16'h1741 : data <= 32'h13017000;
	16'h1742 : data <= 32'h13000000;
	16'h1743 : data <= 32'hb7000080;
	16'h1744 : data <= 32'hb3d12040;
	16'h1745 : data <= 32'h13021200;
	16'h1746 : data <= 32'h93022000;
	16'h1747 : data <= 32'he31452fe;
	16'h1748 : data <= 32'hb70e00ff;
	16'h1749 : data <= 32'h130e7024;
	16'h174a : data <= 32'h6384d101;
	16'h174b : data <= 32'h6f109052;
	16'h174c : data <= 32'h13020000;
	16'h174d : data <= 32'h1301e000;
	16'h174e : data <= 32'h13000000;
	16'h174f : data <= 32'hb7000080;
	16'h1750 : data <= 32'h13000000;
	16'h1751 : data <= 32'hb3d12040;
	16'h1752 : data <= 32'h13021200;
	16'h1753 : data <= 32'h93022000;
	16'h1754 : data <= 32'he31252fe;
	16'h1755 : data <= 32'hb70efeff;
	16'h1756 : data <= 32'h130e8024;
	16'h1757 : data <= 32'h6384d101;
	16'h1758 : data <= 32'h6f10504f;
	16'h1759 : data <= 32'h13020000;
	16'h175a : data <= 32'h1301f001;
	16'h175b : data <= 32'h13000000;
	16'h175c : data <= 32'h13000000;
	16'h175d : data <= 32'hb7000080;
	16'h175e : data <= 32'hb3d12040;
	16'h175f : data <= 32'h13021200;
	16'h1760 : data <= 32'h93022000;
	16'h1761 : data <= 32'he31252fe;
	16'h1762 : data <= 32'h930ef0ff;
	16'h1763 : data <= 32'h130e9024;
	16'h1764 : data <= 32'h6384d101;
	16'h1765 : data <= 32'h6f10104c;
	16'h1766 : data <= 32'h9300f000;
	16'h1767 : data <= 32'h33511040;
	16'h1768 : data <= 32'h930e0000;
	16'h1769 : data <= 32'h130ea024;
	16'h176a : data <= 32'h6304d101;
	16'h176b : data <= 32'h6f10904a;
	16'h176c : data <= 32'h93000002;
	16'h176d : data <= 32'h33d10040;
	16'h176e : data <= 32'h930e0002;
	16'h176f : data <= 32'h130eb024;
	16'h1770 : data <= 32'h6304d101;
	16'h1771 : data <= 32'h6f101049;
	16'h1772 : data <= 32'hb3500040;
	16'h1773 : data <= 32'h930e0000;
	16'h1774 : data <= 32'h130ec024;
	16'h1775 : data <= 32'h6384d001;
	16'h1776 : data <= 32'h6f10d047;
	16'h1777 : data <= 32'h93000040;
	16'h1778 : data <= 32'h37110000;
	16'h1779 : data <= 32'h13010180;
	16'h177a : data <= 32'h33d02040;
	16'h177b : data <= 32'h930e0000;
	16'h177c : data <= 32'h130ed024;
	16'h177d : data <= 32'h6304d001;
	16'h177e : data <= 32'h6f10d045;
	16'h177f : data <= 32'h93000000;
	16'h1780 : data <= 32'h93d10040;
	16'h1781 : data <= 32'h930e0000;
	16'h1782 : data <= 32'h130ee024;
	16'h1783 : data <= 32'h6384d101;
	16'h1784 : data <= 32'h6f105044;
	16'h1785 : data <= 32'hb7000080;
	16'h1786 : data <= 32'h93d11040;
	16'h1787 : data <= 32'hb70e00c0;
	16'h1788 : data <= 32'h130ef024;
	16'h1789 : data <= 32'h6384d101;
	16'h178a : data <= 32'h6f10d042;
	16'h178b : data <= 32'hb7000080;
	16'h178c : data <= 32'h93d17040;
	16'h178d : data <= 32'hb70e00ff;
	16'h178e : data <= 32'h130e0025;
	16'h178f : data <= 32'h6384d101;
	16'h1790 : data <= 32'h6f105041;
	16'h1791 : data <= 32'hb7000080;
	16'h1792 : data <= 32'h93d1e040;
	16'h1793 : data <= 32'hb70efeff;
	16'h1794 : data <= 32'h130e1025;
	16'h1795 : data <= 32'h6384d101;
	16'h1796 : data <= 32'h6f10d03f;
	16'h1797 : data <= 32'hb7000080;
	16'h1798 : data <= 32'h93801000;
	16'h1799 : data <= 32'h93d1f041;
	16'h179a : data <= 32'h930ef0ff;
	16'h179b : data <= 32'h130e2025;
	16'h179c : data <= 32'h6384d101;
	16'h179d : data <= 32'h6f10103e;
	16'h179e : data <= 32'hb7000080;
	16'h179f : data <= 32'h9380f0ff;
	16'h17a0 : data <= 32'h93d10040;
	16'h17a1 : data <= 32'hb70e0080;
	16'h17a2 : data <= 32'h938efeff;
	16'h17a3 : data <= 32'h130e3025;
	16'h17a4 : data <= 32'h6384d101;
	16'h17a5 : data <= 32'h6f10103c;
	16'h17a6 : data <= 32'hb7000080;
	16'h17a7 : data <= 32'h9380f0ff;
	16'h17a8 : data <= 32'h93d11040;
	16'h17a9 : data <= 32'hb70e0040;
	16'h17aa : data <= 32'h938efeff;
	16'h17ab : data <= 32'h130e4025;
	16'h17ac : data <= 32'h6384d101;
	16'h17ad : data <= 32'h6f10103a;
	16'h17ae : data <= 32'hb7000080;
	16'h17af : data <= 32'h9380f0ff;
	16'h17b0 : data <= 32'h93d17040;
	16'h17b1 : data <= 32'hb70e0001;
	16'h17b2 : data <= 32'h938efeff;
	16'h17b3 : data <= 32'h130e5025;
	16'h17b4 : data <= 32'h6384d101;
	16'h17b5 : data <= 32'h6f101038;
	16'h17b6 : data <= 32'hb7000080;
	16'h17b7 : data <= 32'h9380f0ff;
	16'h17b8 : data <= 32'h93d1e040;
	16'h17b9 : data <= 32'hb70e0200;
	16'h17ba : data <= 32'h938efeff;
	16'h17bb : data <= 32'h130e6025;
	16'h17bc : data <= 32'h6384d101;
	16'h17bd : data <= 32'h6f101036;
	16'h17be : data <= 32'hb7000080;
	16'h17bf : data <= 32'h9380f0ff;
	16'h17c0 : data <= 32'h93d1f041;
	16'h17c1 : data <= 32'h930e0000;
	16'h17c2 : data <= 32'h130e7025;
	16'h17c3 : data <= 32'h6384d101;
	16'h17c4 : data <= 32'h6f105034;
	16'h17c5 : data <= 32'hb7808181;
	16'h17c6 : data <= 32'h93801018;
	16'h17c7 : data <= 32'h93d10040;
	16'h17c8 : data <= 32'hb78e8181;
	16'h17c9 : data <= 32'h938e1e18;
	16'h17ca : data <= 32'h130e8025;
	16'h17cb : data <= 32'h6384d101;
	16'h17cc : data <= 32'h6f105032;
	16'h17cd : data <= 32'hb7808181;
	16'h17ce : data <= 32'h93801018;
	16'h17cf : data <= 32'h93d11040;
	16'h17d0 : data <= 32'hb7cec0c0;
	16'h17d1 : data <= 32'h938e0e0c;
	16'h17d2 : data <= 32'h130e9025;
	16'h17d3 : data <= 32'h6384d101;
	16'h17d4 : data <= 32'h6f105030;
	16'h17d5 : data <= 32'hb7808181;
	16'h17d6 : data <= 32'h93801018;
	16'h17d7 : data <= 32'h93d17040;
	16'h17d8 : data <= 32'hb70e03ff;
	16'h17d9 : data <= 32'h938e3e30;
	16'h17da : data <= 32'h130ea025;
	16'h17db : data <= 32'h6384d101;
	16'h17dc : data <= 32'h6f10502e;
	16'h17dd : data <= 32'hb7808181;
	16'h17de : data <= 32'h93801018;
	16'h17df : data <= 32'h93d1e040;
	16'h17e0 : data <= 32'hb70efeff;
	16'h17e1 : data <= 32'h938e6e60;
	16'h17e2 : data <= 32'h130eb025;
	16'h17e3 : data <= 32'h6384d101;
	16'h17e4 : data <= 32'h6f10502c;
	16'h17e5 : data <= 32'hb7808181;
	16'h17e6 : data <= 32'h93801018;
	16'h17e7 : data <= 32'h93d1f041;
	16'h17e8 : data <= 32'h930ef0ff;
	16'h17e9 : data <= 32'h130ec025;
	16'h17ea : data <= 32'h6384d101;
	16'h17eb : data <= 32'h6f10902a;
	16'h17ec : data <= 32'hb7000080;
	16'h17ed : data <= 32'h93d07040;
	16'h17ee : data <= 32'hb70e00ff;
	16'h17ef : data <= 32'h130ed025;
	16'h17f0 : data <= 32'h6384d001;
	16'h17f1 : data <= 32'h6f101029;
	16'h17f2 : data <= 32'h13020000;
	16'h17f3 : data <= 32'hb7000080;
	16'h17f4 : data <= 32'h93d17040;
	16'h17f5 : data <= 32'h13830100;
	16'h17f6 : data <= 32'h13021200;
	16'h17f7 : data <= 32'h93022000;
	16'h17f8 : data <= 32'he31652fe;
	16'h17f9 : data <= 32'hb70e00ff;
	16'h17fa : data <= 32'h130ee025;
	16'h17fb : data <= 32'h6304d301;
	16'h17fc : data <= 32'h6f105026;
	16'h17fd : data <= 32'h13020000;
	16'h17fe : data <= 32'hb7000080;
	16'h17ff : data <= 32'h93d1e040;
	16'h1800 : data <= 32'h13000000;
	16'h1801 : data <= 32'h13830100;
	16'h1802 : data <= 32'h13021200;
	16'h1803 : data <= 32'h93022000;
	16'h1804 : data <= 32'he31452fe;
	16'h1805 : data <= 32'hb70efeff;
	16'h1806 : data <= 32'h130ef025;
	16'h1807 : data <= 32'h6304d301;
	16'h1808 : data <= 32'h6f105023;
	16'h1809 : data <= 32'h13020000;
	16'h180a : data <= 32'hb7000080;
	16'h180b : data <= 32'h93801000;
	16'h180c : data <= 32'h93d1f041;
	16'h180d : data <= 32'h13000000;
	16'h180e : data <= 32'h13000000;
	16'h180f : data <= 32'h13830100;
	16'h1810 : data <= 32'h13021200;
	16'h1811 : data <= 32'h93022000;
	16'h1812 : data <= 32'he31052fe;
	16'h1813 : data <= 32'h930ef0ff;
	16'h1814 : data <= 32'h130e0026;
	16'h1815 : data <= 32'h6304d301;
	16'h1816 : data <= 32'h6f10d01f;
	16'h1817 : data <= 32'h13020000;
	16'h1818 : data <= 32'hb7000080;
	16'h1819 : data <= 32'h93d17040;
	16'h181a : data <= 32'h13021200;
	16'h181b : data <= 32'h93022000;
	16'h181c : data <= 32'he31852fe;
	16'h181d : data <= 32'hb70e00ff;
	16'h181e : data <= 32'h130e1026;
	16'h181f : data <= 32'h6384d101;
	16'h1820 : data <= 32'h6f10501d;
	16'h1821 : data <= 32'h13020000;
	16'h1822 : data <= 32'hb7000080;
	16'h1823 : data <= 32'h13000000;
	16'h1824 : data <= 32'h93d1e040;
	16'h1825 : data <= 32'h13021200;
	16'h1826 : data <= 32'h93022000;
	16'h1827 : data <= 32'he31652fe;
	16'h1828 : data <= 32'hb70efeff;
	16'h1829 : data <= 32'h130e2026;
	16'h182a : data <= 32'h6384d101;
	16'h182b : data <= 32'h6f10901a;
	16'h182c : data <= 32'h13020000;
	16'h182d : data <= 32'hb7000080;
	16'h182e : data <= 32'h93801000;
	16'h182f : data <= 32'h13000000;
	16'h1830 : data <= 32'h13000000;
	16'h1831 : data <= 32'h93d1f041;
	16'h1832 : data <= 32'h13021200;
	16'h1833 : data <= 32'h93022000;
	16'h1834 : data <= 32'he31252fe;
	16'h1835 : data <= 32'h930ef0ff;
	16'h1836 : data <= 32'h130e3026;
	16'h1837 : data <= 32'h6384d101;
	16'h1838 : data <= 32'h6f105017;
	16'h1839 : data <= 32'h9350f041;
	16'h183a : data <= 32'h930e0000;
	16'h183b : data <= 32'h130e4026;
	16'h183c : data <= 32'h6384d001;
	16'h183d : data <= 32'h6f101016;
	16'h183e : data <= 32'h93001002;
	16'h183f : data <= 32'h13d04041;
	16'h1840 : data <= 32'h930e0000;
	16'h1841 : data <= 32'h130e5026;
	16'h1842 : data <= 32'h6304d001;
	16'h1843 : data <= 32'h6f109014;
	16'h1844 : data <= 32'hb780ffff;
	16'h1845 : data <= 32'h13010000;
	16'h1846 : data <= 32'hb3d12000;
	16'h1847 : data <= 32'hb78effff;
	16'h1848 : data <= 32'h130e6026;
	16'h1849 : data <= 32'h6384d101;
	16'h184a : data <= 32'h6f10d012;
	16'h184b : data <= 32'hb780ffff;
	16'h184c : data <= 32'h13011000;
	16'h184d : data <= 32'hb3d12000;
	16'h184e : data <= 32'hb7ceff7f;
	16'h184f : data <= 32'h130e7026;
	16'h1850 : data <= 32'h6384d101;
	16'h1851 : data <= 32'h6f101011;
	16'h1852 : data <= 32'hb780ffff;
	16'h1853 : data <= 32'h13017000;
	16'h1854 : data <= 32'hb3d12000;
	16'h1855 : data <= 32'hb70e0002;
	16'h1856 : data <= 32'h938e0ef0;
	16'h1857 : data <= 32'h130e8026;
	16'h1858 : data <= 32'h6384d101;
	16'h1859 : data <= 32'h6f10100f;
	16'h185a : data <= 32'hb780ffff;
	16'h185b : data <= 32'h1301e000;
	16'h185c : data <= 32'hb3d12000;
	16'h185d : data <= 32'hb70e0400;
	16'h185e : data <= 32'h938eeeff;
	16'h185f : data <= 32'h130e9026;
	16'h1860 : data <= 32'h6384d101;
	16'h1861 : data <= 32'h6f10100d;
	16'h1862 : data <= 32'hb780ffff;
	16'h1863 : data <= 32'h93801000;
	16'h1864 : data <= 32'h1301f000;
	16'h1865 : data <= 32'hb3d12000;
	16'h1866 : data <= 32'hb70e0200;
	16'h1867 : data <= 32'h938efeff;
	16'h1868 : data <= 32'h130ea026;
	16'h1869 : data <= 32'h6384d101;
	16'h186a : data <= 32'h6f10d00a;
	16'h186b : data <= 32'h9300f0ff;
	16'h186c : data <= 32'h13010000;
	16'h186d : data <= 32'hb3d12000;
	16'h186e : data <= 32'h930ef0ff;
	16'h186f : data <= 32'h130eb026;
	16'h1870 : data <= 32'h6384d101;
	16'h1871 : data <= 32'h6f101009;
	16'h1872 : data <= 32'h9300f0ff;
	16'h1873 : data <= 32'h13011000;
	16'h1874 : data <= 32'hb3d12000;
	16'h1875 : data <= 32'hb70e0080;
	16'h1876 : data <= 32'h938efeff;
	16'h1877 : data <= 32'h130ec026;
	16'h1878 : data <= 32'h6384d101;
	16'h1879 : data <= 32'h6f101007;
	16'h187a : data <= 32'h9300f0ff;
	16'h187b : data <= 32'h13017000;
	16'h187c : data <= 32'hb3d12000;
	16'h187d : data <= 32'hb70e0002;
	16'h187e : data <= 32'h938efeff;
	16'h187f : data <= 32'h130ed026;
	16'h1880 : data <= 32'h6384d101;
	16'h1881 : data <= 32'h6f101005;
	16'h1882 : data <= 32'h9300f0ff;
	16'h1883 : data <= 32'h1301e000;
	16'h1884 : data <= 32'hb3d12000;
	16'h1885 : data <= 32'hb70e0400;
	16'h1886 : data <= 32'h938efeff;
	16'h1887 : data <= 32'h130ee026;
	16'h1888 : data <= 32'h6384d101;
	16'h1889 : data <= 32'h6f101003;
	16'h188a : data <= 32'h9300f0ff;
	16'h188b : data <= 32'h1301f001;
	16'h188c : data <= 32'hb3d12000;
	16'h188d : data <= 32'h930e1000;
	16'h188e : data <= 32'h130ef026;
	16'h188f : data <= 32'h6384d101;
	16'h1890 : data <= 32'h6f105001;
	16'h1891 : data <= 32'hb7202121;
	16'h1892 : data <= 32'h93801012;
	16'h1893 : data <= 32'h13010000;
	16'h1894 : data <= 32'hb3d12000;
	16'h1895 : data <= 32'hb72e2121;
	16'h1896 : data <= 32'h938e1e12;
	16'h1897 : data <= 32'h130e0027;
	16'h1898 : data <= 32'h6384d101;
	16'h1899 : data <= 32'h6f10007f;
	16'h189a : data <= 32'hb7202121;
	16'h189b : data <= 32'h93801012;
	16'h189c : data <= 32'h13011000;
	16'h189d : data <= 32'hb3d12000;
	16'h189e : data <= 32'hb79e9010;
	16'h189f : data <= 32'h938e0e09;
	16'h18a0 : data <= 32'h130e1027;
	16'h18a1 : data <= 32'h6384d101;
	16'h18a2 : data <= 32'h6f10c07c;
	16'h18a3 : data <= 32'hb7202121;
	16'h18a4 : data <= 32'h93801012;
	16'h18a5 : data <= 32'h13017000;
	16'h18a6 : data <= 32'hb3d12000;
	16'h18a7 : data <= 32'hb74e4200;
	16'h18a8 : data <= 32'h938e2e24;
	16'h18a9 : data <= 32'h130e2027;
	16'h18aa : data <= 32'h6384d101;
	16'h18ab : data <= 32'h6f10807a;
	16'h18ac : data <= 32'hb7202121;
	16'h18ad : data <= 32'h93801012;
	16'h18ae : data <= 32'h1301e000;
	16'h18af : data <= 32'hb3d12000;
	16'h18b0 : data <= 32'hb78e0000;
	16'h18b1 : data <= 32'h938e4e48;
	16'h18b2 : data <= 32'h130e3027;
	16'h18b3 : data <= 32'h6384d101;
	16'h18b4 : data <= 32'h6f104078;
	16'h18b5 : data <= 32'hb7202121;
	16'h18b6 : data <= 32'h93801012;
	16'h18b7 : data <= 32'h1301f001;
	16'h18b8 : data <= 32'hb3d12000;
	16'h18b9 : data <= 32'h930e0000;
	16'h18ba : data <= 32'h130e4027;
	16'h18bb : data <= 32'h6384d101;
	16'h18bc : data <= 32'h6f104076;
	16'h18bd : data <= 32'hb7202121;
	16'h18be : data <= 32'h93801012;
	16'h18bf : data <= 32'h130100fe;
	16'h18c0 : data <= 32'hb3d12000;
	16'h18c1 : data <= 32'hb72e2121;
	16'h18c2 : data <= 32'h938e1e12;
	16'h18c3 : data <= 32'h130e5027;
	16'h18c4 : data <= 32'h6384d101;
	16'h18c5 : data <= 32'h6f100074;
	16'h18c6 : data <= 32'hb7202121;
	16'h18c7 : data <= 32'h93801012;
	16'h18c8 : data <= 32'h130110fe;
	16'h18c9 : data <= 32'hb3d12000;
	16'h18ca : data <= 32'hb79e9010;
	16'h18cb : data <= 32'h938e0e09;
	16'h18cc : data <= 32'h130e6027;
	16'h18cd : data <= 32'h6384d101;
	16'h18ce : data <= 32'h6f10c071;
	16'h18cf : data <= 32'hb7202121;
	16'h18d0 : data <= 32'h93801012;
	16'h18d1 : data <= 32'h130170fe;
	16'h18d2 : data <= 32'hb3d12000;
	16'h18d3 : data <= 32'hb74e4200;
	16'h18d4 : data <= 32'h938e2e24;
	16'h18d5 : data <= 32'h130e7027;
	16'h18d6 : data <= 32'h6384d101;
	16'h18d7 : data <= 32'h6f10806f;
	16'h18d8 : data <= 32'hb7202121;
	16'h18d9 : data <= 32'h93801012;
	16'h18da : data <= 32'h1301e0fe;
	16'h18db : data <= 32'hb3d12000;
	16'h18dc : data <= 32'hb78e0000;
	16'h18dd : data <= 32'h938e4e48;
	16'h18de : data <= 32'h130e8027;
	16'h18df : data <= 32'h6384d101;
	16'h18e0 : data <= 32'h6f10406d;
	16'h18e1 : data <= 32'hb7202121;
	16'h18e2 : data <= 32'h93801012;
	16'h18e3 : data <= 32'h1301f0ff;
	16'h18e4 : data <= 32'hb3d12000;
	16'h18e5 : data <= 32'h930e0000;
	16'h18e6 : data <= 32'h130e9027;
	16'h18e7 : data <= 32'h6384d101;
	16'h18e8 : data <= 32'h6f10406b;
	16'h18e9 : data <= 32'hb780ffff;
	16'h18ea : data <= 32'h13011000;
	16'h18eb : data <= 32'hb3d02000;
	16'h18ec : data <= 32'hb7ceff7f;
	16'h18ed : data <= 32'h130ea027;
	16'h18ee : data <= 32'h6384d001;
	16'h18ef : data <= 32'h6f108069;
	16'h18f0 : data <= 32'hb780ffff;
	16'h18f1 : data <= 32'h1301e000;
	16'h18f2 : data <= 32'h33d12000;
	16'h18f3 : data <= 32'hb70e0400;
	16'h18f4 : data <= 32'h938eeeff;
	16'h18f5 : data <= 32'h130eb027;
	16'h18f6 : data <= 32'h6304d101;
	16'h18f7 : data <= 32'h6f108067;
	16'h18f8 : data <= 32'h93007000;
	16'h18f9 : data <= 32'hb3d01000;
	16'h18fa : data <= 32'h930e0000;
	16'h18fb : data <= 32'h130ec027;
	16'h18fc : data <= 32'h6384d001;
	16'h18fd : data <= 32'h6f100066;
	16'h18fe : data <= 32'h13020000;
	16'h18ff : data <= 32'hb780ffff;
	16'h1900 : data <= 32'h13011000;
	16'h1901 : data <= 32'hb3d12000;
	16'h1902 : data <= 32'h13830100;
	16'h1903 : data <= 32'h13021200;
	16'h1904 : data <= 32'h93022000;
	16'h1905 : data <= 32'he31452fe;
	16'h1906 : data <= 32'hb7ceff7f;
	16'h1907 : data <= 32'h130ed027;
	16'h1908 : data <= 32'h6304d301;
	16'h1909 : data <= 32'h6f100063;
	16'h190a : data <= 32'h13020000;
	16'h190b : data <= 32'hb780ffff;
	16'h190c : data <= 32'h1301e000;
	16'h190d : data <= 32'hb3d12000;
	16'h190e : data <= 32'h13000000;
	16'h190f : data <= 32'h13830100;
	16'h1910 : data <= 32'h13021200;
	16'h1911 : data <= 32'h93022000;
	16'h1912 : data <= 32'he31252fe;
	16'h1913 : data <= 32'hb70e0400;
	16'h1914 : data <= 32'h938eeeff;
	16'h1915 : data <= 32'h130ee027;
	16'h1916 : data <= 32'h6304d301;
	16'h1917 : data <= 32'h6f10805f;
	16'h1918 : data <= 32'h13020000;
	16'h1919 : data <= 32'hb780ffff;
	16'h191a : data <= 32'h1301f000;
	16'h191b : data <= 32'hb3d12000;
	16'h191c : data <= 32'h13000000;
	16'h191d : data <= 32'h13000000;
	16'h191e : data <= 32'h13830100;
	16'h191f : data <= 32'h13021200;
	16'h1920 : data <= 32'h93022000;
	16'h1921 : data <= 32'he31052fe;
	16'h1922 : data <= 32'hb70e0200;
	16'h1923 : data <= 32'h938efeff;
	16'h1924 : data <= 32'h130ef027;
	16'h1925 : data <= 32'h6304d301;
	16'h1926 : data <= 32'h6f10c05b;
	16'h1927 : data <= 32'h13020000;
	16'h1928 : data <= 32'hb780ffff;
	16'h1929 : data <= 32'h13011000;
	16'h192a : data <= 32'hb3d12000;
	16'h192b : data <= 32'h13021200;
	16'h192c : data <= 32'h93022000;
	16'h192d : data <= 32'he31652fe;
	16'h192e : data <= 32'hb7ceff7f;
	16'h192f : data <= 32'h130e0028;
	16'h1930 : data <= 32'h6384d101;
	16'h1931 : data <= 32'h6f100059;
	16'h1932 : data <= 32'h13020000;
	16'h1933 : data <= 32'hb780ffff;
	16'h1934 : data <= 32'h13017000;
	16'h1935 : data <= 32'h13000000;
	16'h1936 : data <= 32'hb3d12000;
	16'h1937 : data <= 32'h13021200;
	16'h1938 : data <= 32'h93022000;
	16'h1939 : data <= 32'he31452fe;
	16'h193a : data <= 32'hb70e0002;
	16'h193b : data <= 32'h938e0ef0;
	16'h193c : data <= 32'h130e1028;
	16'h193d : data <= 32'h6384d101;
	16'h193e : data <= 32'h6f10c055;
	16'h193f : data <= 32'h13020000;
	16'h1940 : data <= 32'hb780ffff;
	16'h1941 : data <= 32'h1301f000;
	16'h1942 : data <= 32'h13000000;
	16'h1943 : data <= 32'h13000000;
	16'h1944 : data <= 32'hb3d12000;
	16'h1945 : data <= 32'h13021200;
	16'h1946 : data <= 32'h93022000;
	16'h1947 : data <= 32'he31252fe;
	16'h1948 : data <= 32'hb70e0200;
	16'h1949 : data <= 32'h938efeff;
	16'h194a : data <= 32'h130e2028;
	16'h194b : data <= 32'h6384d101;
	16'h194c : data <= 32'h6f104052;
	16'h194d : data <= 32'h13020000;
	16'h194e : data <= 32'hb780ffff;
	16'h194f : data <= 32'h13000000;
	16'h1950 : data <= 32'h13011000;
	16'h1951 : data <= 32'hb3d12000;
	16'h1952 : data <= 32'h13021200;
	16'h1953 : data <= 32'h93022000;
	16'h1954 : data <= 32'he31452fe;
	16'h1955 : data <= 32'hb7ceff7f;
	16'h1956 : data <= 32'h130e3028;
	16'h1957 : data <= 32'h6384d101;
	16'h1958 : data <= 32'h6f10404f;
	16'h1959 : data <= 32'h13020000;
	16'h195a : data <= 32'hb780ffff;
	16'h195b : data <= 32'h13000000;
	16'h195c : data <= 32'h13017000;
	16'h195d : data <= 32'h13000000;
	16'h195e : data <= 32'hb3d12000;
	16'h195f : data <= 32'h13021200;
	16'h1960 : data <= 32'h93022000;
	16'h1961 : data <= 32'he31252fe;
	16'h1962 : data <= 32'hb70e0002;
	16'h1963 : data <= 32'h938e0ef0;
	16'h1964 : data <= 32'h130e4028;
	16'h1965 : data <= 32'h6384d101;
	16'h1966 : data <= 32'h6f10c04b;
	16'h1967 : data <= 32'h13020000;
	16'h1968 : data <= 32'hb780ffff;
	16'h1969 : data <= 32'h13000000;
	16'h196a : data <= 32'h13000000;
	16'h196b : data <= 32'h1301f000;
	16'h196c : data <= 32'hb3d12000;
	16'h196d : data <= 32'h13021200;
	16'h196e : data <= 32'h93022000;
	16'h196f : data <= 32'he31252fe;
	16'h1970 : data <= 32'hb70e0200;
	16'h1971 : data <= 32'h938efeff;
	16'h1972 : data <= 32'h130e5028;
	16'h1973 : data <= 32'h6384d101;
	16'h1974 : data <= 32'h6f104048;
	16'h1975 : data <= 32'h13020000;
	16'h1976 : data <= 32'h13011000;
	16'h1977 : data <= 32'hb780ffff;
	16'h1978 : data <= 32'hb3d12000;
	16'h1979 : data <= 32'h13021200;
	16'h197a : data <= 32'h93022000;
	16'h197b : data <= 32'he31652fe;
	16'h197c : data <= 32'hb7ceff7f;
	16'h197d : data <= 32'h130e6028;
	16'h197e : data <= 32'h6384d101;
	16'h197f : data <= 32'h6f108045;
	16'h1980 : data <= 32'h13020000;
	16'h1981 : data <= 32'h13017000;
	16'h1982 : data <= 32'hb780ffff;
	16'h1983 : data <= 32'h13000000;
	16'h1984 : data <= 32'hb3d12000;
	16'h1985 : data <= 32'h13021200;
	16'h1986 : data <= 32'h93022000;
	16'h1987 : data <= 32'he31452fe;
	16'h1988 : data <= 32'hb70e0002;
	16'h1989 : data <= 32'h938e0ef0;
	16'h198a : data <= 32'h130e7028;
	16'h198b : data <= 32'h6384d101;
	16'h198c : data <= 32'h6f104042;
	16'h198d : data <= 32'h13020000;
	16'h198e : data <= 32'h1301f000;
	16'h198f : data <= 32'hb780ffff;
	16'h1990 : data <= 32'h13000000;
	16'h1991 : data <= 32'h13000000;
	16'h1992 : data <= 32'hb3d12000;
	16'h1993 : data <= 32'h13021200;
	16'h1994 : data <= 32'h93022000;
	16'h1995 : data <= 32'he31252fe;
	16'h1996 : data <= 32'hb70e0200;
	16'h1997 : data <= 32'h938efeff;
	16'h1998 : data <= 32'h130e8028;
	16'h1999 : data <= 32'h6384d101;
	16'h199a : data <= 32'h6f10c03e;
	16'h199b : data <= 32'h13020000;
	16'h199c : data <= 32'h13011000;
	16'h199d : data <= 32'h13000000;
	16'h199e : data <= 32'hb780ffff;
	16'h199f : data <= 32'hb3d12000;
	16'h19a0 : data <= 32'h13021200;
	16'h19a1 : data <= 32'h93022000;
	16'h19a2 : data <= 32'he31452fe;
	16'h19a3 : data <= 32'hb7ceff7f;
	16'h19a4 : data <= 32'h130e9028;
	16'h19a5 : data <= 32'h6384d101;
	16'h19a6 : data <= 32'h6f10c03b;
	16'h19a7 : data <= 32'h13020000;
	16'h19a8 : data <= 32'h13017000;
	16'h19a9 : data <= 32'h13000000;
	16'h19aa : data <= 32'hb780ffff;
	16'h19ab : data <= 32'h13000000;
	16'h19ac : data <= 32'hb3d12000;
	16'h19ad : data <= 32'h13021200;
	16'h19ae : data <= 32'h93022000;
	16'h19af : data <= 32'he31252fe;
	16'h19b0 : data <= 32'hb70e0002;
	16'h19b1 : data <= 32'h938e0ef0;
	16'h19b2 : data <= 32'h130ea028;
	16'h19b3 : data <= 32'h6384d101;
	16'h19b4 : data <= 32'h6f104038;
	16'h19b5 : data <= 32'h13020000;
	16'h19b6 : data <= 32'h1301f000;
	16'h19b7 : data <= 32'h13000000;
	16'h19b8 : data <= 32'h13000000;
	16'h19b9 : data <= 32'hb780ffff;
	16'h19ba : data <= 32'hb3d12000;
	16'h19bb : data <= 32'h13021200;
	16'h19bc : data <= 32'h93022000;
	16'h19bd : data <= 32'he31252fe;
	16'h19be : data <= 32'hb70e0200;
	16'h19bf : data <= 32'h938efeff;
	16'h19c0 : data <= 32'h130eb028;
	16'h19c1 : data <= 32'h6384d101;
	16'h19c2 : data <= 32'h6f10c034;
	16'h19c3 : data <= 32'h9300f000;
	16'h19c4 : data <= 32'h33511000;
	16'h19c5 : data <= 32'h930e0000;
	16'h19c6 : data <= 32'h130ec028;
	16'h19c7 : data <= 32'h6304d101;
	16'h19c8 : data <= 32'h6f104033;
	16'h19c9 : data <= 32'h93000002;
	16'h19ca : data <= 32'h33d10000;
	16'h19cb : data <= 32'h930e0002;
	16'h19cc : data <= 32'h130ed028;
	16'h19cd : data <= 32'h6304d101;
	16'h19ce : data <= 32'h6f10c031;
	16'h19cf : data <= 32'hb3500000;
	16'h19d0 : data <= 32'h930e0000;
	16'h19d1 : data <= 32'h130ee028;
	16'h19d2 : data <= 32'h6384d001;
	16'h19d3 : data <= 32'h6f108030;
	16'h19d4 : data <= 32'h93000040;
	16'h19d5 : data <= 32'h37110000;
	16'h19d6 : data <= 32'h13010180;
	16'h19d7 : data <= 32'h33d02000;
	16'h19d8 : data <= 32'h930e0000;
	16'h19d9 : data <= 32'h130ef028;
	16'h19da : data <= 32'h6304d001;
	16'h19db : data <= 32'h6f10802e;
	16'h19dc : data <= 32'hb780ffff;
	16'h19dd : data <= 32'h93d10000;
	16'h19de : data <= 32'hb78effff;
	16'h19df : data <= 32'h130e0029;
	16'h19e0 : data <= 32'h6384d101;
	16'h19e1 : data <= 32'h6f10002d;
	16'h19e2 : data <= 32'hb780ffff;
	16'h19e3 : data <= 32'h93d11000;
	16'h19e4 : data <= 32'hb7ceff7f;
	16'h19e5 : data <= 32'h130e1029;
	16'h19e6 : data <= 32'h6384d101;
	16'h19e7 : data <= 32'h6f10802b;
	16'h19e8 : data <= 32'hb780ffff;
	16'h19e9 : data <= 32'h93d17000;
	16'h19ea : data <= 32'hb70e0002;
	16'h19eb : data <= 32'h938e0ef0;
	16'h19ec : data <= 32'h130e2029;
	16'h19ed : data <= 32'h6384d101;
	16'h19ee : data <= 32'h6f10c029;
	16'h19ef : data <= 32'hb780ffff;
	16'h19f0 : data <= 32'h93d1e000;
	16'h19f1 : data <= 32'hb70e0400;
	16'h19f2 : data <= 32'h938eeeff;
	16'h19f3 : data <= 32'h130e3029;
	16'h19f4 : data <= 32'h6384d101;
	16'h19f5 : data <= 32'h6f100028;
	16'h19f6 : data <= 32'hb780ffff;
	16'h19f7 : data <= 32'h93801000;
	16'h19f8 : data <= 32'h93d1f000;
	16'h19f9 : data <= 32'hb70e0200;
	16'h19fa : data <= 32'h938efeff;
	16'h19fb : data <= 32'h130e4029;
	16'h19fc : data <= 32'h6384d101;
	16'h19fd : data <= 32'h6f100026;
	16'h19fe : data <= 32'h9300f0ff;
	16'h19ff : data <= 32'h93d10000;
	16'h1a00 : data <= 32'h930ef0ff;
	16'h1a01 : data <= 32'h130e5029;
	16'h1a02 : data <= 32'h6384d101;
	16'h1a03 : data <= 32'h6f108024;
	16'h1a04 : data <= 32'h9300f0ff;
	16'h1a05 : data <= 32'h93d11000;
	16'h1a06 : data <= 32'hb70e0080;
	16'h1a07 : data <= 32'h938efeff;
	16'h1a08 : data <= 32'h130e6029;
	16'h1a09 : data <= 32'h6384d101;
	16'h1a0a : data <= 32'h6f10c022;
	16'h1a0b : data <= 32'h9300f0ff;
	16'h1a0c : data <= 32'h93d17000;
	16'h1a0d : data <= 32'hb70e0002;
	16'h1a0e : data <= 32'h938efeff;
	16'h1a0f : data <= 32'h130e7029;
	16'h1a10 : data <= 32'h6384d101;
	16'h1a11 : data <= 32'h6f100021;
	16'h1a12 : data <= 32'h9300f0ff;
	16'h1a13 : data <= 32'h93d1e000;
	16'h1a14 : data <= 32'hb70e0400;
	16'h1a15 : data <= 32'h938efeff;
	16'h1a16 : data <= 32'h130e8029;
	16'h1a17 : data <= 32'h6384d101;
	16'h1a18 : data <= 32'h6f10401f;
	16'h1a19 : data <= 32'h9300f0ff;
	16'h1a1a : data <= 32'h93d1f001;
	16'h1a1b : data <= 32'h930e1000;
	16'h1a1c : data <= 32'h130e9029;
	16'h1a1d : data <= 32'h6384d101;
	16'h1a1e : data <= 32'h6f10c01d;
	16'h1a1f : data <= 32'hb7202121;
	16'h1a20 : data <= 32'h93801012;
	16'h1a21 : data <= 32'h93d10000;
	16'h1a22 : data <= 32'hb72e2121;
	16'h1a23 : data <= 32'h938e1e12;
	16'h1a24 : data <= 32'h130ea029;
	16'h1a25 : data <= 32'h6384d101;
	16'h1a26 : data <= 32'h6f10c01b;
	16'h1a27 : data <= 32'hb7202121;
	16'h1a28 : data <= 32'h93801012;
	16'h1a29 : data <= 32'h93d11000;
	16'h1a2a : data <= 32'hb79e9010;
	16'h1a2b : data <= 32'h938e0e09;
	16'h1a2c : data <= 32'h130eb029;
	16'h1a2d : data <= 32'h6384d101;
	16'h1a2e : data <= 32'h6f10c019;
	16'h1a2f : data <= 32'hb7202121;
	16'h1a30 : data <= 32'h93801012;
	16'h1a31 : data <= 32'h93d17000;
	16'h1a32 : data <= 32'hb74e4200;
	16'h1a33 : data <= 32'h938e2e24;
	16'h1a34 : data <= 32'h130ec029;
	16'h1a35 : data <= 32'h6384d101;
	16'h1a36 : data <= 32'h6f10c017;
	16'h1a37 : data <= 32'hb7202121;
	16'h1a38 : data <= 32'h93801012;
	16'h1a39 : data <= 32'h93d1e000;
	16'h1a3a : data <= 32'hb78e0000;
	16'h1a3b : data <= 32'h938e4e48;
	16'h1a3c : data <= 32'h130ed029;
	16'h1a3d : data <= 32'h6384d101;
	16'h1a3e : data <= 32'h6f10c015;
	16'h1a3f : data <= 32'hb7202121;
	16'h1a40 : data <= 32'h93801012;
	16'h1a41 : data <= 32'h93d1f001;
	16'h1a42 : data <= 32'h930e0000;
	16'h1a43 : data <= 32'h130ee029;
	16'h1a44 : data <= 32'h6384d101;
	16'h1a45 : data <= 32'h6f100014;
	16'h1a46 : data <= 32'hb780ffff;
	16'h1a47 : data <= 32'h93d01000;
	16'h1a48 : data <= 32'hb7ceff7f;
	16'h1a49 : data <= 32'h130ef029;
	16'h1a4a : data <= 32'h6384d001;
	16'h1a4b : data <= 32'h6f108012;
	16'h1a4c : data <= 32'h13020000;
	16'h1a4d : data <= 32'hb780ffff;
	16'h1a4e : data <= 32'h93d11000;
	16'h1a4f : data <= 32'h13830100;
	16'h1a50 : data <= 32'h13021200;
	16'h1a51 : data <= 32'h93022000;
	16'h1a52 : data <= 32'he31652fe;
	16'h1a53 : data <= 32'hb7ceff7f;
	16'h1a54 : data <= 32'h130e002a;
	16'h1a55 : data <= 32'h6304d301;
	16'h1a56 : data <= 32'h6f10c00f;
	16'h1a57 : data <= 32'h13020000;
	16'h1a58 : data <= 32'hb780ffff;
	16'h1a59 : data <= 32'h93d1e000;
	16'h1a5a : data <= 32'h13000000;
	16'h1a5b : data <= 32'h13830100;
	16'h1a5c : data <= 32'h13021200;
	16'h1a5d : data <= 32'h93022000;
	16'h1a5e : data <= 32'he31452fe;
	16'h1a5f : data <= 32'hb70e0400;
	16'h1a60 : data <= 32'h938eeeff;
	16'h1a61 : data <= 32'h130e102a;
	16'h1a62 : data <= 32'h6304d301;
	16'h1a63 : data <= 32'h6f10800c;
	16'h1a64 : data <= 32'h13020000;
	16'h1a65 : data <= 32'hb780ffff;
	16'h1a66 : data <= 32'h93d1f000;
	16'h1a67 : data <= 32'h13000000;
	16'h1a68 : data <= 32'h13000000;
	16'h1a69 : data <= 32'h13830100;
	16'h1a6a : data <= 32'h13021200;
	16'h1a6b : data <= 32'h93022000;
	16'h1a6c : data <= 32'he31252fe;
	16'h1a6d : data <= 32'hb70e0200;
	16'h1a6e : data <= 32'h938efeff;
	16'h1a6f : data <= 32'h130e202a;
	16'h1a70 : data <= 32'h6304d301;
	16'h1a71 : data <= 32'h6f100009;
	16'h1a72 : data <= 32'h13020000;
	16'h1a73 : data <= 32'hb780ffff;
	16'h1a74 : data <= 32'h93d11000;
	16'h1a75 : data <= 32'h13021200;
	16'h1a76 : data <= 32'h93022000;
	16'h1a77 : data <= 32'he31852fe;
	16'h1a78 : data <= 32'hb7ceff7f;
	16'h1a79 : data <= 32'h130e302a;
	16'h1a7a : data <= 32'h6384d101;
	16'h1a7b : data <= 32'h6f108006;
	16'h1a7c : data <= 32'h13020000;
	16'h1a7d : data <= 32'hb780ffff;
	16'h1a7e : data <= 32'h13000000;
	16'h1a7f : data <= 32'h93d1e000;
	16'h1a80 : data <= 32'h13021200;
	16'h1a81 : data <= 32'h93022000;
	16'h1a82 : data <= 32'he31652fe;
	16'h1a83 : data <= 32'hb70e0400;
	16'h1a84 : data <= 32'h938eeeff;
	16'h1a85 : data <= 32'h130e402a;
	16'h1a86 : data <= 32'h6384d101;
	16'h1a87 : data <= 32'h6f108003;
	16'h1a88 : data <= 32'h13020000;
	16'h1a89 : data <= 32'hb780ffff;
	16'h1a8a : data <= 32'h13000000;
	16'h1a8b : data <= 32'h13000000;
	16'h1a8c : data <= 32'h93d1f000;
	16'h1a8d : data <= 32'h13021200;
	16'h1a8e : data <= 32'h93022000;
	16'h1a8f : data <= 32'he31452fe;
	16'h1a90 : data <= 32'hb70e0200;
	16'h1a91 : data <= 32'h938efeff;
	16'h1a92 : data <= 32'h130e502a;
	16'h1a93 : data <= 32'h6384d101;
	16'h1a94 : data <= 32'h6f104000;
	16'h1a95 : data <= 32'h9350f001;
	16'h1a96 : data <= 32'h930e0000;
	16'h1a97 : data <= 32'h130e602a;
	16'h1a98 : data <= 32'he39ad07f;
	16'h1a99 : data <= 32'h93001002;
	16'h1a9a : data <= 32'h13d04001;
	16'h1a9b : data <= 32'h930e0000;
	16'h1a9c : data <= 32'h130e702a;
	16'h1a9d : data <= 32'he310d07f;
	16'h1a9e : data <= 32'h93000000;
	16'h1a9f : data <= 32'h13010000;
	16'h1aa0 : data <= 32'hb3812040;
	16'h1aa1 : data <= 32'h930e0000;
	16'h1aa2 : data <= 32'h130e802a;
	16'h1aa3 : data <= 32'he394d17d;
	16'h1aa4 : data <= 32'h93001000;
	16'h1aa5 : data <= 32'h13011000;
	16'h1aa6 : data <= 32'hb3812040;
	16'h1aa7 : data <= 32'h930e0000;
	16'h1aa8 : data <= 32'h130e902a;
	16'h1aa9 : data <= 32'he398d17b;
	16'h1aaa : data <= 32'h93003000;
	16'h1aab : data <= 32'h13017000;
	16'h1aac : data <= 32'hb3812040;
	16'h1aad : data <= 32'h930ec0ff;
	16'h1aae : data <= 32'h130ea02a;
	16'h1aaf : data <= 32'he39cd179;
	16'h1ab0 : data <= 32'h93000000;
	16'h1ab1 : data <= 32'h3781ffff;
	16'h1ab2 : data <= 32'hb3812040;
	16'h1ab3 : data <= 32'hb78e0000;
	16'h1ab4 : data <= 32'h130eb02a;
	16'h1ab5 : data <= 32'he390d179;
	16'h1ab6 : data <= 32'hb7000080;
	16'h1ab7 : data <= 32'h13010000;
	16'h1ab8 : data <= 32'hb3812040;
	16'h1ab9 : data <= 32'hb70e0080;
	16'h1aba : data <= 32'h130ec02a;
	16'h1abb : data <= 32'he394d177;
	16'h1abc : data <= 32'hb7000080;
	16'h1abd : data <= 32'h3781ffff;
	16'h1abe : data <= 32'hb3812040;
	16'h1abf : data <= 32'hb78e0080;
	16'h1ac0 : data <= 32'h130ed02a;
	16'h1ac1 : data <= 32'he398d175;
	16'h1ac2 : data <= 32'h93000000;
	16'h1ac3 : data <= 32'h37810000;
	16'h1ac4 : data <= 32'h1301f1ff;
	16'h1ac5 : data <= 32'hb3812040;
	16'h1ac6 : data <= 32'hb78effff;
	16'h1ac7 : data <= 32'h938e1e00;
	16'h1ac8 : data <= 32'h130ee02a;
	16'h1ac9 : data <= 32'he398d173;
	16'h1aca : data <= 32'hb7000080;
	16'h1acb : data <= 32'h9380f0ff;
	16'h1acc : data <= 32'h13010000;
	16'h1acd : data <= 32'hb3812040;
	16'h1ace : data <= 32'hb70e0080;
	16'h1acf : data <= 32'h938efeff;
	16'h1ad0 : data <= 32'h130ef02a;
	16'h1ad1 : data <= 32'he398d171;
	16'h1ad2 : data <= 32'hb7000080;
	16'h1ad3 : data <= 32'h9380f0ff;
	16'h1ad4 : data <= 32'h37810000;
	16'h1ad5 : data <= 32'h1301f1ff;
	16'h1ad6 : data <= 32'hb3812040;
	16'h1ad7 : data <= 32'hb78eff7f;
	16'h1ad8 : data <= 32'h130e002b;
	16'h1ad9 : data <= 32'he398d16f;
	16'h1ada : data <= 32'hb7000080;
	16'h1adb : data <= 32'h37810000;
	16'h1adc : data <= 32'h1301f1ff;
	16'h1add : data <= 32'hb3812040;
	16'h1ade : data <= 32'hb78eff7f;
	16'h1adf : data <= 32'h938e1e00;
	16'h1ae0 : data <= 32'h130e102b;
	16'h1ae1 : data <= 32'he398d16d;
	16'h1ae2 : data <= 32'hb7000080;
	16'h1ae3 : data <= 32'h9380f0ff;
	16'h1ae4 : data <= 32'h3781ffff;
	16'h1ae5 : data <= 32'hb3812040;
	16'h1ae6 : data <= 32'hb78e0080;
	16'h1ae7 : data <= 32'h938efeff;
	16'h1ae8 : data <= 32'h130e202b;
	16'h1ae9 : data <= 32'he398d16b;
	16'h1aea : data <= 32'h93000000;
	16'h1aeb : data <= 32'h1301f0ff;
	16'h1aec : data <= 32'hb3812040;
	16'h1aed : data <= 32'h930e1000;
	16'h1aee : data <= 32'h130e302b;
	16'h1aef : data <= 32'he39cd169;
	16'h1af0 : data <= 32'h9300f0ff;
	16'h1af1 : data <= 32'h13011000;
	16'h1af2 : data <= 32'hb3812040;
	16'h1af3 : data <= 32'h930ee0ff;
	16'h1af4 : data <= 32'h130e402b;
	16'h1af5 : data <= 32'he390d169;
	16'h1af6 : data <= 32'h9300f0ff;
	16'h1af7 : data <= 32'h1301f0ff;
	16'h1af8 : data <= 32'hb3812040;
	16'h1af9 : data <= 32'h930e0000;
	16'h1afa : data <= 32'h130e502b;
	16'h1afb : data <= 32'he394d167;
	16'h1afc : data <= 32'h9300d000;
	16'h1afd : data <= 32'h1301b000;
	16'h1afe : data <= 32'hb3802040;
	16'h1aff : data <= 32'h930e2000;
	16'h1b00 : data <= 32'h130e602b;
	16'h1b01 : data <= 32'he398d065;
	16'h1b02 : data <= 32'h9300e000;
	16'h1b03 : data <= 32'h1301b000;
	16'h1b04 : data <= 32'h33812040;
	16'h1b05 : data <= 32'h930e3000;
	16'h1b06 : data <= 32'h130e702b;
	16'h1b07 : data <= 32'he31cd163;
	16'h1b08 : data <= 32'h9300d000;
	16'h1b09 : data <= 32'hb3801040;
	16'h1b0a : data <= 32'h930e0000;
	16'h1b0b : data <= 32'h130e802b;
	16'h1b0c : data <= 32'he392d063;
	16'h1b0d : data <= 32'h13020000;
	16'h1b0e : data <= 32'h9300d000;
	16'h1b0f : data <= 32'h1301b000;
	16'h1b10 : data <= 32'hb3812040;
	16'h1b11 : data <= 32'h13830100;
	16'h1b12 : data <= 32'h13021200;
	16'h1b13 : data <= 32'h93022000;
	16'h1b14 : data <= 32'he31452fe;
	16'h1b15 : data <= 32'h930e2000;
	16'h1b16 : data <= 32'h130e902b;
	16'h1b17 : data <= 32'he31cd35f;
	16'h1b18 : data <= 32'h13020000;
	16'h1b19 : data <= 32'h9300e000;
	16'h1b1a : data <= 32'h1301b000;
	16'h1b1b : data <= 32'hb3812040;
	16'h1b1c : data <= 32'h13000000;
	16'h1b1d : data <= 32'h13830100;
	16'h1b1e : data <= 32'h13021200;
	16'h1b1f : data <= 32'h93022000;
	16'h1b20 : data <= 32'he31252fe;
	16'h1b21 : data <= 32'h930e3000;
	16'h1b22 : data <= 32'h130ea02b;
	16'h1b23 : data <= 32'he314d35d;
	16'h1b24 : data <= 32'h13020000;
	16'h1b25 : data <= 32'h9300f000;
	16'h1b26 : data <= 32'h1301b000;
	16'h1b27 : data <= 32'hb3812040;
	16'h1b28 : data <= 32'h13000000;
	16'h1b29 : data <= 32'h13000000;
	16'h1b2a : data <= 32'h13830100;
	16'h1b2b : data <= 32'h13021200;
	16'h1b2c : data <= 32'h93022000;
	16'h1b2d : data <= 32'he31052fe;
	16'h1b2e : data <= 32'h930e4000;
	16'h1b2f : data <= 32'h130eb02b;
	16'h1b30 : data <= 32'he31ad359;
	16'h1b31 : data <= 32'h13020000;
	16'h1b32 : data <= 32'h9300d000;
	16'h1b33 : data <= 32'h1301b000;
	16'h1b34 : data <= 32'hb3812040;
	16'h1b35 : data <= 32'h13021200;
	16'h1b36 : data <= 32'h93022000;
	16'h1b37 : data <= 32'he31652fe;
	16'h1b38 : data <= 32'h930e2000;
	16'h1b39 : data <= 32'h130ec02b;
	16'h1b3a : data <= 32'he396d157;
	16'h1b3b : data <= 32'h13020000;
	16'h1b3c : data <= 32'h9300e000;
	16'h1b3d : data <= 32'h1301b000;
	16'h1b3e : data <= 32'h13000000;
	16'h1b3f : data <= 32'hb3812040;
	16'h1b40 : data <= 32'h13021200;
	16'h1b41 : data <= 32'h93022000;
	16'h1b42 : data <= 32'he31452fe;
	16'h1b43 : data <= 32'h930e3000;
	16'h1b44 : data <= 32'h130ed02b;
	16'h1b45 : data <= 32'he390d155;
	16'h1b46 : data <= 32'h13020000;
	16'h1b47 : data <= 32'h9300f000;
	16'h1b48 : data <= 32'h1301b000;
	16'h1b49 : data <= 32'h13000000;
	16'h1b4a : data <= 32'h13000000;
	16'h1b4b : data <= 32'hb3812040;
	16'h1b4c : data <= 32'h13021200;
	16'h1b4d : data <= 32'h93022000;
	16'h1b4e : data <= 32'he31252fe;
	16'h1b4f : data <= 32'h930e4000;
	16'h1b50 : data <= 32'h130ee02b;
	16'h1b51 : data <= 32'he398d151;
	16'h1b52 : data <= 32'h13020000;
	16'h1b53 : data <= 32'h9300d000;
	16'h1b54 : data <= 32'h13000000;
	16'h1b55 : data <= 32'h1301b000;
	16'h1b56 : data <= 32'hb3812040;
	16'h1b57 : data <= 32'h13021200;
	16'h1b58 : data <= 32'h93022000;
	16'h1b59 : data <= 32'he31452fe;
	16'h1b5a : data <= 32'h930e2000;
	16'h1b5b : data <= 32'h130ef02b;
	16'h1b5c : data <= 32'he392d14f;
	16'h1b5d : data <= 32'h13020000;
	16'h1b5e : data <= 32'h9300e000;
	16'h1b5f : data <= 32'h13000000;
	16'h1b60 : data <= 32'h1301b000;
	16'h1b61 : data <= 32'h13000000;
	16'h1b62 : data <= 32'hb3812040;
	16'h1b63 : data <= 32'h13021200;
	16'h1b64 : data <= 32'h93022000;
	16'h1b65 : data <= 32'he31252fe;
	16'h1b66 : data <= 32'h930e3000;
	16'h1b67 : data <= 32'h130e002c;
	16'h1b68 : data <= 32'he39ad14b;
	16'h1b69 : data <= 32'h13020000;
	16'h1b6a : data <= 32'h9300f000;
	16'h1b6b : data <= 32'h13000000;
	16'h1b6c : data <= 32'h13000000;
	16'h1b6d : data <= 32'h1301b000;
	16'h1b6e : data <= 32'hb3812040;
	16'h1b6f : data <= 32'h13021200;
	16'h1b70 : data <= 32'h93022000;
	16'h1b71 : data <= 32'he31252fe;
	16'h1b72 : data <= 32'h930e4000;
	16'h1b73 : data <= 32'h130e102c;
	16'h1b74 : data <= 32'he392d149;
	16'h1b75 : data <= 32'h13020000;
	16'h1b76 : data <= 32'h1301b000;
	16'h1b77 : data <= 32'h9300d000;
	16'h1b78 : data <= 32'hb3812040;
	16'h1b79 : data <= 32'h13021200;
	16'h1b7a : data <= 32'h93022000;
	16'h1b7b : data <= 32'he31652fe;
	16'h1b7c : data <= 32'h930e2000;
	16'h1b7d : data <= 32'h130e202c;
	16'h1b7e : data <= 32'he39ed145;
	16'h1b7f : data <= 32'h13020000;
	16'h1b80 : data <= 32'h1301b000;
	16'h1b81 : data <= 32'h9300e000;
	16'h1b82 : data <= 32'h13000000;
	16'h1b83 : data <= 32'hb3812040;
	16'h1b84 : data <= 32'h13021200;
	16'h1b85 : data <= 32'h93022000;
	16'h1b86 : data <= 32'he31452fe;
	16'h1b87 : data <= 32'h930e3000;
	16'h1b88 : data <= 32'h130e302c;
	16'h1b89 : data <= 32'he398d143;
	16'h1b8a : data <= 32'h13020000;
	16'h1b8b : data <= 32'h1301b000;
	16'h1b8c : data <= 32'h9300f000;
	16'h1b8d : data <= 32'h13000000;
	16'h1b8e : data <= 32'h13000000;
	16'h1b8f : data <= 32'hb3812040;
	16'h1b90 : data <= 32'h13021200;
	16'h1b91 : data <= 32'h93022000;
	16'h1b92 : data <= 32'he31252fe;
	16'h1b93 : data <= 32'h930e4000;
	16'h1b94 : data <= 32'h130e402c;
	16'h1b95 : data <= 32'he390d141;
	16'h1b96 : data <= 32'h13020000;
	16'h1b97 : data <= 32'h1301b000;
	16'h1b98 : data <= 32'h13000000;
	16'h1b99 : data <= 32'h9300d000;
	16'h1b9a : data <= 32'hb3812040;
	16'h1b9b : data <= 32'h13021200;
	16'h1b9c : data <= 32'h93022000;
	16'h1b9d : data <= 32'he31452fe;
	16'h1b9e : data <= 32'h930e2000;
	16'h1b9f : data <= 32'h130e502c;
	16'h1ba0 : data <= 32'he39ad13d;
	16'h1ba1 : data <= 32'h13020000;
	16'h1ba2 : data <= 32'h1301b000;
	16'h1ba3 : data <= 32'h13000000;
	16'h1ba4 : data <= 32'h9300e000;
	16'h1ba5 : data <= 32'h13000000;
	16'h1ba6 : data <= 32'hb3812040;
	16'h1ba7 : data <= 32'h13021200;
	16'h1ba8 : data <= 32'h93022000;
	16'h1ba9 : data <= 32'he31252fe;
	16'h1baa : data <= 32'h930e3000;
	16'h1bab : data <= 32'h130e602c;
	16'h1bac : data <= 32'he392d13b;
	16'h1bad : data <= 32'h13020000;
	16'h1bae : data <= 32'h1301b000;
	16'h1baf : data <= 32'h13000000;
	16'h1bb0 : data <= 32'h13000000;
	16'h1bb1 : data <= 32'h9300f000;
	16'h1bb2 : data <= 32'hb3812040;
	16'h1bb3 : data <= 32'h13021200;
	16'h1bb4 : data <= 32'h93022000;
	16'h1bb5 : data <= 32'he31252fe;
	16'h1bb6 : data <= 32'h930e4000;
	16'h1bb7 : data <= 32'h130e702c;
	16'h1bb8 : data <= 32'he39ad137;
	16'h1bb9 : data <= 32'h930010ff;
	16'h1bba : data <= 32'h33011040;
	16'h1bbb : data <= 32'h930ef000;
	16'h1bbc : data <= 32'h130e802c;
	16'h1bbd : data <= 32'he310d137;
	16'h1bbe : data <= 32'h93000002;
	16'h1bbf : data <= 32'h33810040;
	16'h1bc0 : data <= 32'h930e0002;
	16'h1bc1 : data <= 32'h130e902c;
	16'h1bc2 : data <= 32'he316d135;
	16'h1bc3 : data <= 32'hb3000040;
	16'h1bc4 : data <= 32'h930e0000;
	16'h1bc5 : data <= 32'h130ea02c;
	16'h1bc6 : data <= 32'he39ed033;
	16'h1bc7 : data <= 32'h93000001;
	16'h1bc8 : data <= 32'h1301e001;
	16'h1bc9 : data <= 32'h33802040;
	16'h1bca : data <= 32'h930e0000;
	16'h1bcb : data <= 32'h130eb02c;
	16'h1bcc : data <= 32'he312d033;
	16'h1bcd : data <= 32'h97100000;
	16'h1bce : data <= 32'h93802011;
	16'h1bcf : data <= 32'h3701aa00;
	16'h1bd0 : data <= 32'h1301a10a;
	16'h1bd1 : data <= 32'h23a02000;
	16'h1bd2 : data <= 32'h83a10000;
	16'h1bd3 : data <= 32'hb70eaa00;
	16'h1bd4 : data <= 32'h938eae0a;
	16'h1bd5 : data <= 32'h130ec02c;
	16'h1bd6 : data <= 32'he39ed12f;
	16'h1bd7 : data <= 32'h97100000;
	16'h1bd8 : data <= 32'h9380a00e;
	16'h1bd9 : data <= 32'h37b100aa;
	16'h1bda : data <= 32'h130101a0;
	16'h1bdb : data <= 32'h23a22000;
	16'h1bdc : data <= 32'h83a14000;
	16'h1bdd : data <= 32'hb7be00aa;
	16'h1bde : data <= 32'h938e0ea0;
	16'h1bdf : data <= 32'h130ed02c;
	16'h1be0 : data <= 32'he39ad12d;
	16'h1be1 : data <= 32'h97100000;
	16'h1be2 : data <= 32'h9380200c;
	16'h1be3 : data <= 32'h3711a00a;
	16'h1be4 : data <= 32'h130101aa;
	16'h1be5 : data <= 32'h23a42000;
	16'h1be6 : data <= 32'h83a18000;
	16'h1be7 : data <= 32'hb71ea00a;
	16'h1be8 : data <= 32'h938e0eaa;
	16'h1be9 : data <= 32'h130ee02c;
	16'h1bea : data <= 32'he396d12b;
	16'h1beb : data <= 32'h97100000;
	16'h1bec : data <= 32'h9380a009;
	16'h1bed : data <= 32'h37a10aa0;
	16'h1bee : data <= 32'h1301a100;
	16'h1bef : data <= 32'h23a62000;
	16'h1bf0 : data <= 32'h83a1c000;
	16'h1bf1 : data <= 32'hb7ae0aa0;
	16'h1bf2 : data <= 32'h938eae00;
	16'h1bf3 : data <= 32'h130ef02c;
	16'h1bf4 : data <= 32'he392d129;
	16'h1bf5 : data <= 32'h97100000;
	16'h1bf6 : data <= 32'h9380e008;
	16'h1bf7 : data <= 32'h3701aa00;
	16'h1bf8 : data <= 32'h1301a10a;
	16'h1bf9 : data <= 32'h23aa20fe;
	16'h1bfa : data <= 32'h83a140ff;
	16'h1bfb : data <= 32'hb70eaa00;
	16'h1bfc : data <= 32'h938eae0a;
	16'h1bfd : data <= 32'h130e002d;
	16'h1bfe : data <= 32'he39ed125;
	16'h1bff : data <= 32'h97100000;
	16'h1c00 : data <= 32'h93806006;
	16'h1c01 : data <= 32'h37b100aa;
	16'h1c02 : data <= 32'h130101a0;
	16'h1c03 : data <= 32'h23ac20fe;
	16'h1c04 : data <= 32'h83a180ff;
	16'h1c05 : data <= 32'hb7be00aa;
	16'h1c06 : data <= 32'h938e0ea0;
	16'h1c07 : data <= 32'h130e102d;
	16'h1c08 : data <= 32'he39ad123;
	16'h1c09 : data <= 32'h97100000;
	16'h1c0a : data <= 32'h9380e003;
	16'h1c0b : data <= 32'h3711a00a;
	16'h1c0c : data <= 32'h130101aa;
	16'h1c0d : data <= 32'h23ae20fe;
	16'h1c0e : data <= 32'h83a1c0ff;
	16'h1c0f : data <= 32'hb71ea00a;
	16'h1c10 : data <= 32'h938e0eaa;
	16'h1c11 : data <= 32'h130e202d;
	16'h1c12 : data <= 32'he396d121;
	16'h1c13 : data <= 32'h97100000;
	16'h1c14 : data <= 32'h93806001;
	16'h1c15 : data <= 32'h37a10aa0;
	16'h1c16 : data <= 32'h1301a100;
	16'h1c17 : data <= 32'h23a02000;
	16'h1c18 : data <= 32'h83a10000;
	16'h1c19 : data <= 32'hb7ae0aa0;
	16'h1c1a : data <= 32'h938eae00;
	16'h1c1b : data <= 32'h130e302d;
	16'h1c1c : data <= 32'he392d11f;
	16'h1c1d : data <= 32'h97100000;
	16'h1c1e : data <= 32'h938020ff;
	16'h1c1f : data <= 32'h37513412;
	16'h1c20 : data <= 32'h13018167;
	16'h1c21 : data <= 32'h138200fe;
	16'h1c22 : data <= 32'h23202202;
	16'h1c23 : data <= 32'h83a10000;
	16'h1c24 : data <= 32'hb75e3412;
	16'h1c25 : data <= 32'h938e8e67;
	16'h1c26 : data <= 32'h130e402d;
	16'h1c27 : data <= 32'he39cd11b;
	16'h1c28 : data <= 32'h97100000;
	16'h1c29 : data <= 32'h938060fc;
	16'h1c2a : data <= 32'h37312158;
	16'h1c2b : data <= 32'h13018109;
	16'h1c2c : data <= 32'h9380d0ff;
	16'h1c2d : data <= 32'ha3a32000;
	16'h1c2e : data <= 32'h17120000;
	16'h1c2f : data <= 32'h130222fb;
	16'h1c30 : data <= 32'h83210200;
	16'h1c31 : data <= 32'hb73e2158;
	16'h1c32 : data <= 32'h938e8e09;
	16'h1c33 : data <= 32'h130e502d;
	16'h1c34 : data <= 32'he392d119;
	16'h1c35 : data <= 32'h130e602d;
	16'h1c36 : data <= 32'h13020000;
	16'h1c37 : data <= 32'hb7d0bbaa;
	16'h1c38 : data <= 32'h9380d0cd;
	16'h1c39 : data <= 32'h17110000;
	16'h1c3a : data <= 32'h130121f6;
	16'h1c3b : data <= 32'h23201100;
	16'h1c3c : data <= 32'h83210100;
	16'h1c3d : data <= 32'hb7debbaa;
	16'h1c3e : data <= 32'h938edecd;
	16'h1c3f : data <= 32'he39cd115;
	16'h1c40 : data <= 32'h13021200;
	16'h1c41 : data <= 32'h93022000;
	16'h1c42 : data <= 32'he31a52fc;
	16'h1c43 : data <= 32'h130e702d;
	16'h1c44 : data <= 32'h13020000;
	16'h1c45 : data <= 32'hb7c0abda;
	16'h1c46 : data <= 32'h9380d0cc;
	16'h1c47 : data <= 32'h17110000;
	16'h1c48 : data <= 32'h1301a1f2;
	16'h1c49 : data <= 32'h13000000;
	16'h1c4a : data <= 32'h23221100;
	16'h1c4b : data <= 32'h83214100;
	16'h1c4c : data <= 32'hb7ceabda;
	16'h1c4d : data <= 32'h938edecc;
	16'h1c4e : data <= 32'he39ed111;
	16'h1c4f : data <= 32'h13021200;
	16'h1c50 : data <= 32'h93022000;
	16'h1c51 : data <= 32'he31852fc;
	16'h1c52 : data <= 32'h130e802d;
	16'h1c53 : data <= 32'h13020000;
	16'h1c54 : data <= 32'hb7c0aadd;
	16'h1c55 : data <= 32'h9380c0bc;
	16'h1c56 : data <= 32'h17110000;
	16'h1c57 : data <= 32'h1301e1ee;
	16'h1c58 : data <= 32'h13000000;
	16'h1c59 : data <= 32'h13000000;
	16'h1c5a : data <= 32'h23241100;
	16'h1c5b : data <= 32'h83218100;
	16'h1c5c : data <= 32'hb7ceaadd;
	16'h1c5d : data <= 32'h938ecebc;
	16'h1c5e : data <= 32'he39ed10d;
	16'h1c5f : data <= 32'h13021200;
	16'h1c60 : data <= 32'h93022000;
	16'h1c61 : data <= 32'he31652fc;
	16'h1c62 : data <= 32'h130e902d;
	16'h1c63 : data <= 32'h13020000;
	16'h1c64 : data <= 32'hb7b0dacd;
	16'h1c65 : data <= 32'h9380c0bb;
	16'h1c66 : data <= 32'h13000000;
	16'h1c67 : data <= 32'h17110000;
	16'h1c68 : data <= 32'h1301a1ea;
	16'h1c69 : data <= 32'h23261100;
	16'h1c6a : data <= 32'h8321c100;
	16'h1c6b : data <= 32'hb7bedacd;
	16'h1c6c : data <= 32'h938ecebb;
	16'h1c6d : data <= 32'he390d10b;
	16'h1c6e : data <= 32'h13021200;
	16'h1c6f : data <= 32'h93022000;
	16'h1c70 : data <= 32'he31852fc;
	16'h1c71 : data <= 32'h130ea02d;
	16'h1c72 : data <= 32'h13020000;
	16'h1c73 : data <= 32'hb7b0ddcc;
	16'h1c74 : data <= 32'h9380b0ab;
	16'h1c75 : data <= 32'h13000000;
	16'h1c76 : data <= 32'h17110000;
	16'h1c77 : data <= 32'h1301e1e6;
	16'h1c78 : data <= 32'h13000000;
	16'h1c79 : data <= 32'h23281100;
	16'h1c7a : data <= 32'h83210101;
	16'h1c7b : data <= 32'hb7beddcc;
	16'h1c7c : data <= 32'h938ebeab;
	16'h1c7d : data <= 32'he390d107;
	16'h1c7e : data <= 32'h13021200;
	16'h1c7f : data <= 32'h93022000;
	16'h1c80 : data <= 32'he31652fc;
	16'h1c81 : data <= 32'h130eb02d;
	16'h1c82 : data <= 32'h13020000;
	16'h1c83 : data <= 32'hb7e0cdbc;
	16'h1c84 : data <= 32'h9380b0aa;
	16'h1c85 : data <= 32'h13000000;
	16'h1c86 : data <= 32'h13000000;
	16'h1c87 : data <= 32'h17110000;
	16'h1c88 : data <= 32'h1301a1e2;
	16'h1c89 : data <= 32'h232a1100;
	16'h1c8a : data <= 32'h83214101;
	16'h1c8b : data <= 32'hb7eecdbc;
	16'h1c8c : data <= 32'h938ebeaa;
	16'h1c8d : data <= 32'he390d103;
	16'h1c8e : data <= 32'h13021200;
	16'h1c8f : data <= 32'h93022000;
	16'h1c90 : data <= 32'he31652fc;
	16'h1c91 : data <= 32'h130ec02d;
	16'h1c92 : data <= 32'h13020000;
	16'h1c93 : data <= 32'h17110000;
	16'h1c94 : data <= 32'h1301a1df;
	16'h1c95 : data <= 32'hb7201100;
	16'h1c96 : data <= 32'h93803023;
	16'h1c97 : data <= 32'h23201100;
	16'h1c98 : data <= 32'h83210100;
	16'h1c99 : data <= 32'hb72e1100;
	16'h1c9a : data <= 32'h938e3e23;
	16'h1c9b : data <= 32'h6394d17f;
	16'h1c9c : data <= 32'h13021200;
	16'h1c9d : data <= 32'h93022000;
	16'h1c9e : data <= 32'he31a52fc;
	16'h1c9f : data <= 32'h130ed02d;
	16'h1ca0 : data <= 32'h13020000;
	16'h1ca1 : data <= 32'h17110000;
	16'h1ca2 : data <= 32'h130121dc;
	16'h1ca3 : data <= 32'hb7100130;
	16'h1ca4 : data <= 32'h93803022;
	16'h1ca5 : data <= 32'h13000000;
	16'h1ca6 : data <= 32'h23221100;
	16'h1ca7 : data <= 32'h83214100;
	16'h1ca8 : data <= 32'hb71e0130;
	16'h1ca9 : data <= 32'h938e3e22;
	16'h1caa : data <= 32'h6396d17b;
	16'h1cab : data <= 32'h13021200;
	16'h1cac : data <= 32'h93022000;
	16'h1cad : data <= 32'he31852fc;
	16'h1cae : data <= 32'h130ee02d;
	16'h1caf : data <= 32'h13020000;
	16'h1cb0 : data <= 32'h17110000;
	16'h1cb1 : data <= 32'h130161d8;
	16'h1cb2 : data <= 32'hb7100033;
	16'h1cb3 : data <= 32'h93802012;
	16'h1cb4 : data <= 32'h13000000;
	16'h1cb5 : data <= 32'h13000000;
	16'h1cb6 : data <= 32'h23241100;
	16'h1cb7 : data <= 32'h83218100;
	16'h1cb8 : data <= 32'hb71e0033;
	16'h1cb9 : data <= 32'h938e2e12;
	16'h1cba : data <= 32'h6396d177;
	16'h1cbb : data <= 32'h13021200;
	16'h1cbc : data <= 32'h93022000;
	16'h1cbd : data <= 32'he31652fc;
	16'h1cbe : data <= 32'h130ef02d;
	16'h1cbf : data <= 32'h13020000;
	16'h1cc0 : data <= 32'h17110000;
	16'h1cc1 : data <= 32'h130161d4;
	16'h1cc2 : data <= 32'h13000000;
	16'h1cc3 : data <= 32'hb7003023;
	16'h1cc4 : data <= 32'h93802011;
	16'h1cc5 : data <= 32'h23261100;
	16'h1cc6 : data <= 32'h8321c100;
	16'h1cc7 : data <= 32'hb70e3023;
	16'h1cc8 : data <= 32'h938e2e11;
	16'h1cc9 : data <= 32'h6398d173;
	16'h1cca : data <= 32'h13021200;
	16'h1ccb : data <= 32'h93022000;
	16'h1ccc : data <= 32'he31852fc;
	16'h1ccd : data <= 32'h130e002e;
	16'h1cce : data <= 32'h13020000;
	16'h1ccf : data <= 32'h17110000;
	16'h1cd0 : data <= 32'h1301a1d0;
	16'h1cd1 : data <= 32'h13000000;
	16'h1cd2 : data <= 32'hb7003322;
	16'h1cd3 : data <= 32'h93801001;
	16'h1cd4 : data <= 32'h13000000;
	16'h1cd5 : data <= 32'h23281100;
	16'h1cd6 : data <= 32'h83210101;
	16'h1cd7 : data <= 32'hb70e3322;
	16'h1cd8 : data <= 32'h938e1e01;
	16'h1cd9 : data <= 32'h6398d16f;
	16'h1cda : data <= 32'h13021200;
	16'h1cdb : data <= 32'h93022000;
	16'h1cdc : data <= 32'he31652fc;
	16'h1cdd : data <= 32'h130e102e;
	16'h1cde : data <= 32'h13020000;
	16'h1cdf : data <= 32'h17110000;
	16'h1ce0 : data <= 32'h1301a1cc;
	16'h1ce1 : data <= 32'h13000000;
	16'h1ce2 : data <= 32'h13000000;
	16'h1ce3 : data <= 32'hb7302312;
	16'h1ce4 : data <= 32'h93801000;
	16'h1ce5 : data <= 32'h232a1100;
	16'h1ce6 : data <= 32'h83214101;
	16'h1ce7 : data <= 32'hb73e2312;
	16'h1ce8 : data <= 32'h938e1e00;
	16'h1ce9 : data <= 32'h6398d16b;
	16'h1cea : data <= 32'h13021200;
	16'h1ceb : data <= 32'h93022000;
	16'h1cec : data <= 32'he31652fc;
	16'h1ced : data <= 32'hb70001ff;
	16'h1cee : data <= 32'h938000f0;
	16'h1cef : data <= 32'h37110f0f;
	16'h1cf0 : data <= 32'h1301f1f0;
	16'h1cf1 : data <= 32'hb3c12000;
	16'h1cf2 : data <= 32'hb7fe0ff0;
	16'h1cf3 : data <= 32'h938efe00;
	16'h1cf4 : data <= 32'h130e202e;
	16'h1cf5 : data <= 32'h6390d169;
	16'h1cf6 : data <= 32'hb710f00f;
	16'h1cf7 : data <= 32'h938000ff;
	16'h1cf8 : data <= 32'h37f1f0f0;
	16'h1cf9 : data <= 32'h1301010f;
	16'h1cfa : data <= 32'hb3c12000;
	16'h1cfb : data <= 32'hb70e01ff;
	16'h1cfc : data <= 32'h938e0ef0;
	16'h1cfd : data <= 32'h130e302e;
	16'h1cfe : data <= 32'h639ed165;
	16'h1cff : data <= 32'hb700ff00;
	16'h1d00 : data <= 32'h9380f00f;
	16'h1d01 : data <= 32'h37110f0f;
	16'h1d02 : data <= 32'h1301f1f0;
	16'h1d03 : data <= 32'hb3c12000;
	16'h1d04 : data <= 32'hb71ef00f;
	16'h1d05 : data <= 32'h938e0eff;
	16'h1d06 : data <= 32'h130e402e;
	16'h1d07 : data <= 32'h639cd163;
	16'h1d08 : data <= 32'hb7f00ff0;
	16'h1d09 : data <= 32'h9380f000;
	16'h1d0a : data <= 32'h37f1f0f0;
	16'h1d0b : data <= 32'h1301010f;
	16'h1d0c : data <= 32'hb3c12000;
	16'h1d0d : data <= 32'hb70eff00;
	16'h1d0e : data <= 32'h938efe0f;
	16'h1d0f : data <= 32'h130e502e;
	16'h1d10 : data <= 32'h639ad161;
	16'h1d11 : data <= 32'hb70001ff;
	16'h1d12 : data <= 32'h938000f0;
	16'h1d13 : data <= 32'h37110f0f;
	16'h1d14 : data <= 32'h1301f1f0;
	16'h1d15 : data <= 32'hb3c02000;
	16'h1d16 : data <= 32'hb7fe0ff0;
	16'h1d17 : data <= 32'h938efe00;
	16'h1d18 : data <= 32'h130e602e;
	16'h1d19 : data <= 32'h6398d05f;
	16'h1d1a : data <= 32'hb70001ff;
	16'h1d1b : data <= 32'h938000f0;
	16'h1d1c : data <= 32'h37110f0f;
	16'h1d1d : data <= 32'h1301f1f0;
	16'h1d1e : data <= 32'h33c12000;
	16'h1d1f : data <= 32'hb7fe0ff0;
	16'h1d20 : data <= 32'h938efe00;
	16'h1d21 : data <= 32'h130e702e;
	16'h1d22 : data <= 32'h6316d15d;
	16'h1d23 : data <= 32'hb70001ff;
	16'h1d24 : data <= 32'h938000f0;
	16'h1d25 : data <= 32'hb3c01000;
	16'h1d26 : data <= 32'h930e0000;
	16'h1d27 : data <= 32'h130e802e;
	16'h1d28 : data <= 32'h639ad05b;
	16'h1d29 : data <= 32'h13020000;
	16'h1d2a : data <= 32'hb70001ff;
	16'h1d2b : data <= 32'h938000f0;
	16'h1d2c : data <= 32'h37110f0f;
	16'h1d2d : data <= 32'h1301f1f0;
	16'h1d2e : data <= 32'hb3c12000;
	16'h1d2f : data <= 32'h13830100;
	16'h1d30 : data <= 32'h13021200;
	16'h1d31 : data <= 32'h93022000;
	16'h1d32 : data <= 32'he31052fe;
	16'h1d33 : data <= 32'hb7fe0ff0;
	16'h1d34 : data <= 32'h938efe00;
	16'h1d35 : data <= 32'h130e902e;
	16'h1d36 : data <= 32'h631ed357;
	16'h1d37 : data <= 32'h13020000;
	16'h1d38 : data <= 32'hb710f00f;
	16'h1d39 : data <= 32'h938000ff;
	16'h1d3a : data <= 32'h37f1f0f0;
	16'h1d3b : data <= 32'h1301010f;
	16'h1d3c : data <= 32'hb3c12000;
	16'h1d3d : data <= 32'h13000000;
	16'h1d3e : data <= 32'h13830100;
	16'h1d3f : data <= 32'h13021200;
	16'h1d40 : data <= 32'h93022000;
	16'h1d41 : data <= 32'he31e52fc;
	16'h1d42 : data <= 32'hb70e01ff;
	16'h1d43 : data <= 32'h938e0ef0;
	16'h1d44 : data <= 32'h130ea02e;
	16'h1d45 : data <= 32'h6310d355;
	16'h1d46 : data <= 32'h13020000;
	16'h1d47 : data <= 32'hb700ff00;
	16'h1d48 : data <= 32'h9380f00f;
	16'h1d49 : data <= 32'h37110f0f;
	16'h1d4a : data <= 32'h1301f1f0;
	16'h1d4b : data <= 32'hb3c12000;
	16'h1d4c : data <= 32'h13000000;
	16'h1d4d : data <= 32'h13000000;
	16'h1d4e : data <= 32'h13830100;
	16'h1d4f : data <= 32'h13021200;
	16'h1d50 : data <= 32'h93022000;
	16'h1d51 : data <= 32'he31c52fc;
	16'h1d52 : data <= 32'hb71ef00f;
	16'h1d53 : data <= 32'h938e0eff;
	16'h1d54 : data <= 32'h130eb02e;
	16'h1d55 : data <= 32'h6310d351;
	16'h1d56 : data <= 32'h13020000;
	16'h1d57 : data <= 32'hb70001ff;
	16'h1d58 : data <= 32'h938000f0;
	16'h1d59 : data <= 32'h37110f0f;
	16'h1d5a : data <= 32'h1301f1f0;
	16'h1d5b : data <= 32'hb3c12000;
	16'h1d5c : data <= 32'h13021200;
	16'h1d5d : data <= 32'h93022000;
	16'h1d5e : data <= 32'he31252fe;
	16'h1d5f : data <= 32'hb7fe0ff0;
	16'h1d60 : data <= 32'h938efe00;
	16'h1d61 : data <= 32'h130ec02e;
	16'h1d62 : data <= 32'h6396d14d;
	16'h1d63 : data <= 32'h13020000;
	16'h1d64 : data <= 32'hb710f00f;
	16'h1d65 : data <= 32'h938000ff;
	16'h1d66 : data <= 32'h37f1f0f0;
	16'h1d67 : data <= 32'h1301010f;
	16'h1d68 : data <= 32'h13000000;
	16'h1d69 : data <= 32'hb3c12000;
	16'h1d6a : data <= 32'h13021200;
	16'h1d6b : data <= 32'h93022000;
	16'h1d6c : data <= 32'he31052fe;
	16'h1d6d : data <= 32'hb70e01ff;
	16'h1d6e : data <= 32'h938e0ef0;
	16'h1d6f : data <= 32'h130ed02e;
	16'h1d70 : data <= 32'h639ad149;
	16'h1d71 : data <= 32'h13020000;
	16'h1d72 : data <= 32'hb700ff00;
	16'h1d73 : data <= 32'h9380f00f;
	16'h1d74 : data <= 32'h37110f0f;
	16'h1d75 : data <= 32'h1301f1f0;
	16'h1d76 : data <= 32'h13000000;
	16'h1d77 : data <= 32'h13000000;
	16'h1d78 : data <= 32'hb3c12000;
	16'h1d79 : data <= 32'h13021200;
	16'h1d7a : data <= 32'h93022000;
	16'h1d7b : data <= 32'he31e52fc;
	16'h1d7c : data <= 32'hb71ef00f;
	16'h1d7d : data <= 32'h938e0eff;
	16'h1d7e : data <= 32'h130ee02e;
	16'h1d7f : data <= 32'h639cd145;
	16'h1d80 : data <= 32'h13020000;
	16'h1d81 : data <= 32'hb70001ff;
	16'h1d82 : data <= 32'h938000f0;
	16'h1d83 : data <= 32'h13000000;
	16'h1d84 : data <= 32'h37110f0f;
	16'h1d85 : data <= 32'h1301f1f0;
	16'h1d86 : data <= 32'hb3c12000;
	16'h1d87 : data <= 32'h13021200;
	16'h1d88 : data <= 32'h93022000;
	16'h1d89 : data <= 32'he31052fe;
	16'h1d8a : data <= 32'hb7fe0ff0;
	16'h1d8b : data <= 32'h938efe00;
	16'h1d8c : data <= 32'h130ef02e;
	16'h1d8d : data <= 32'h6390d143;
	16'h1d8e : data <= 32'h13020000;
	16'h1d8f : data <= 32'hb710f00f;
	16'h1d90 : data <= 32'h938000ff;
	16'h1d91 : data <= 32'h13000000;
	16'h1d92 : data <= 32'h37f1f0f0;
	16'h1d93 : data <= 32'h1301010f;
	16'h1d94 : data <= 32'h13000000;
	16'h1d95 : data <= 32'hb3c12000;
	16'h1d96 : data <= 32'h13021200;
	16'h1d97 : data <= 32'h93022000;
	16'h1d98 : data <= 32'he31e52fc;
	16'h1d99 : data <= 32'hb70e01ff;
	16'h1d9a : data <= 32'h938e0ef0;
	16'h1d9b : data <= 32'h130e002f;
	16'h1d9c : data <= 32'h6392d13f;
	16'h1d9d : data <= 32'h13020000;
	16'h1d9e : data <= 32'hb700ff00;
	16'h1d9f : data <= 32'h9380f00f;
	16'h1da0 : data <= 32'h13000000;
	16'h1da1 : data <= 32'h13000000;
	16'h1da2 : data <= 32'h37110f0f;
	16'h1da3 : data <= 32'h1301f1f0;
	16'h1da4 : data <= 32'hb3c12000;
	16'h1da5 : data <= 32'h13021200;
	16'h1da6 : data <= 32'h93022000;
	16'h1da7 : data <= 32'he31e52fc;
	16'h1da8 : data <= 32'hb71ef00f;
	16'h1da9 : data <= 32'h938e0eff;
	16'h1daa : data <= 32'h130e102f;
	16'h1dab : data <= 32'h6394d13b;
	16'h1dac : data <= 32'h13020000;
	16'h1dad : data <= 32'h37110f0f;
	16'h1dae : data <= 32'h1301f1f0;
	16'h1daf : data <= 32'hb70001ff;
	16'h1db0 : data <= 32'h938000f0;
	16'h1db1 : data <= 32'hb3c12000;
	16'h1db2 : data <= 32'h13021200;
	16'h1db3 : data <= 32'h93022000;
	16'h1db4 : data <= 32'he31252fe;
	16'h1db5 : data <= 32'hb7fe0ff0;
	16'h1db6 : data <= 32'h938efe00;
	16'h1db7 : data <= 32'h130e202f;
	16'h1db8 : data <= 32'h639ad137;
	16'h1db9 : data <= 32'h13020000;
	16'h1dba : data <= 32'h37f1f0f0;
	16'h1dbb : data <= 32'h1301010f;
	16'h1dbc : data <= 32'hb710f00f;
	16'h1dbd : data <= 32'h938000ff;
	16'h1dbe : data <= 32'h13000000;
	16'h1dbf : data <= 32'hb3c12000;
	16'h1dc0 : data <= 32'h13021200;
	16'h1dc1 : data <= 32'h93022000;
	16'h1dc2 : data <= 32'he31052fe;
	16'h1dc3 : data <= 32'hb70e01ff;
	16'h1dc4 : data <= 32'h938e0ef0;
	16'h1dc5 : data <= 32'h130e302f;
	16'h1dc6 : data <= 32'h639ed133;
	16'h1dc7 : data <= 32'h13020000;
	16'h1dc8 : data <= 32'h37110f0f;
	16'h1dc9 : data <= 32'h1301f1f0;
	16'h1dca : data <= 32'hb700ff00;
	16'h1dcb : data <= 32'h9380f00f;
	16'h1dcc : data <= 32'h13000000;
	16'h1dcd : data <= 32'h13000000;
	16'h1dce : data <= 32'hb3c12000;
	16'h1dcf : data <= 32'h13021200;
	16'h1dd0 : data <= 32'h93022000;
	16'h1dd1 : data <= 32'he31e52fc;
	16'h1dd2 : data <= 32'hb71ef00f;
	16'h1dd3 : data <= 32'h938e0eff;
	16'h1dd4 : data <= 32'h130e402f;
	16'h1dd5 : data <= 32'h6390d131;
	16'h1dd6 : data <= 32'h13020000;
	16'h1dd7 : data <= 32'h37110f0f;
	16'h1dd8 : data <= 32'h1301f1f0;
	16'h1dd9 : data <= 32'h13000000;
	16'h1dda : data <= 32'hb70001ff;
	16'h1ddb : data <= 32'h938000f0;
	16'h1ddc : data <= 32'hb3c12000;
	16'h1ddd : data <= 32'h13021200;
	16'h1dde : data <= 32'h93022000;
	16'h1ddf : data <= 32'he31052fe;
	16'h1de0 : data <= 32'hb7fe0ff0;
	16'h1de1 : data <= 32'h938efe00;
	16'h1de2 : data <= 32'h130e502f;
	16'h1de3 : data <= 32'h6394d12d;
	16'h1de4 : data <= 32'h13020000;
	16'h1de5 : data <= 32'h37f1f0f0;
	16'h1de6 : data <= 32'h1301010f;
	16'h1de7 : data <= 32'h13000000;
	16'h1de8 : data <= 32'hb710f00f;
	16'h1de9 : data <= 32'h938000ff;
	16'h1dea : data <= 32'h13000000;
	16'h1deb : data <= 32'hb3c12000;
	16'h1dec : data <= 32'h13021200;
	16'h1ded : data <= 32'h93022000;
	16'h1dee : data <= 32'he31e52fc;
	16'h1def : data <= 32'hb70e01ff;
	16'h1df0 : data <= 32'h938e0ef0;
	16'h1df1 : data <= 32'h130e602f;
	16'h1df2 : data <= 32'h6396d129;
	16'h1df3 : data <= 32'h13020000;
	16'h1df4 : data <= 32'h37110f0f;
	16'h1df5 : data <= 32'h1301f1f0;
	16'h1df6 : data <= 32'h13000000;
	16'h1df7 : data <= 32'h13000000;
	16'h1df8 : data <= 32'hb700ff00;
	16'h1df9 : data <= 32'h9380f00f;
	16'h1dfa : data <= 32'hb3c12000;
	16'h1dfb : data <= 32'h13021200;
	16'h1dfc : data <= 32'h93022000;
	16'h1dfd : data <= 32'he31e52fc;
	16'h1dfe : data <= 32'hb71ef00f;
	16'h1dff : data <= 32'h938e0eff;
	16'h1e00 : data <= 32'h130e702f;
	16'h1e01 : data <= 32'h6398d125;
	16'h1e02 : data <= 32'hb70001ff;
	16'h1e03 : data <= 32'h938000f0;
	16'h1e04 : data <= 32'h33411000;
	16'h1e05 : data <= 32'hb70e01ff;
	16'h1e06 : data <= 32'h938e0ef0;
	16'h1e07 : data <= 32'h130e802f;
	16'h1e08 : data <= 32'h631ad123;
	16'h1e09 : data <= 32'hb700ff00;
	16'h1e0a : data <= 32'h9380f00f;
	16'h1e0b : data <= 32'h33c10000;
	16'h1e0c : data <= 32'hb70eff00;
	16'h1e0d : data <= 32'h938efe0f;
	16'h1e0e : data <= 32'h130e902f;
	16'h1e0f : data <= 32'h631cd121;
	16'h1e10 : data <= 32'hb3400000;
	16'h1e11 : data <= 32'h930e0000;
	16'h1e12 : data <= 32'h130ea02f;
	16'h1e13 : data <= 32'h6394d021;
	16'h1e14 : data <= 32'hb7101111;
	16'h1e15 : data <= 32'h93801011;
	16'h1e16 : data <= 32'h37212222;
	16'h1e17 : data <= 32'h13012122;
	16'h1e18 : data <= 32'h33c02000;
	16'h1e19 : data <= 32'h930e0000;
	16'h1e1a : data <= 32'h130eb02f;
	16'h1e1b : data <= 32'h6314d01f;
	16'h1e1c : data <= 32'hb710ff00;
	16'h1e1d : data <= 32'h938000f0;
	16'h1e1e : data <= 32'h93c1f0f0;
	16'h1e1f : data <= 32'hb7fe00ff;
	16'h1e20 : data <= 32'h938efe00;
	16'h1e21 : data <= 32'h130ec02f;
	16'h1e22 : data <= 32'h6396d11d;
	16'h1e23 : data <= 32'hb710f00f;
	16'h1e24 : data <= 32'h938000ff;
	16'h1e25 : data <= 32'h93c1000f;
	16'h1e26 : data <= 32'hb71ef00f;
	16'h1e27 : data <= 32'h938e0ef0;
	16'h1e28 : data <= 32'h130ed02f;
	16'h1e29 : data <= 32'h6398d11b;
	16'h1e2a : data <= 32'hb710ff00;
	16'h1e2b : data <= 32'h9380f08f;
	16'h1e2c : data <= 32'h93c1f070;
	16'h1e2d : data <= 32'hb71eff00;
	16'h1e2e : data <= 32'h938e0eff;
	16'h1e2f : data <= 32'h130ee02f;
	16'h1e30 : data <= 32'h639ad119;
	16'h1e31 : data <= 32'hb7f00ff0;
	16'h1e32 : data <= 32'h9380f000;
	16'h1e33 : data <= 32'h93c1000f;
	16'h1e34 : data <= 32'hb7fe0ff0;
	16'h1e35 : data <= 32'h938efe0f;
	16'h1e36 : data <= 32'h130ef02f;
	16'h1e37 : data <= 32'h639cd117;
	16'h1e38 : data <= 32'hb7f000ff;
	16'h1e39 : data <= 32'h93800070;
	16'h1e3a : data <= 32'h93c0f070;
	16'h1e3b : data <= 32'hb7fe00ff;
	16'h1e3c : data <= 32'h938efe00;
	16'h1e3d : data <= 32'h130e0030;
	16'h1e3e : data <= 32'h639ed015;
	16'h1e3f : data <= 32'h13020000;
	16'h1e40 : data <= 32'hb710f00f;
	16'h1e41 : data <= 32'h938000ff;
	16'h1e42 : data <= 32'h93c1000f;
	16'h1e43 : data <= 32'h13830100;
	16'h1e44 : data <= 32'h13021200;
	16'h1e45 : data <= 32'h93022000;
	16'h1e46 : data <= 32'he31452fe;
	16'h1e47 : data <= 32'hb71ef00f;
	16'h1e48 : data <= 32'h938e0ef0;
	16'h1e49 : data <= 32'h130e1030;
	16'h1e4a : data <= 32'h6316d313;
	16'h1e4b : data <= 32'h13020000;
	16'h1e4c : data <= 32'hb710ff00;
	16'h1e4d : data <= 32'h9380f08f;
	16'h1e4e : data <= 32'h93c1f070;
	16'h1e4f : data <= 32'h13000000;
	16'h1e50 : data <= 32'h13830100;
	16'h1e51 : data <= 32'h13021200;
	16'h1e52 : data <= 32'h93022000;
	16'h1e53 : data <= 32'he31252fe;
	16'h1e54 : data <= 32'hb71eff00;
	16'h1e55 : data <= 32'h938e0eff;
	16'h1e56 : data <= 32'h130e2030;
	16'h1e57 : data <= 32'h631cd30f;
	16'h1e58 : data <= 32'h13020000;
	16'h1e59 : data <= 32'hb7f00ff0;
	16'h1e5a : data <= 32'h9380f000;
	16'h1e5b : data <= 32'h93c1000f;
	16'h1e5c : data <= 32'h13000000;
	16'h1e5d : data <= 32'h13000000;
	16'h1e5e : data <= 32'h13830100;
	16'h1e5f : data <= 32'h13021200;
	16'h1e60 : data <= 32'h93022000;
	16'h1e61 : data <= 32'he31052fe;
	16'h1e62 : data <= 32'hb7fe0ff0;
	16'h1e63 : data <= 32'h938efe0f;
	16'h1e64 : data <= 32'h130e3030;
	16'h1e65 : data <= 32'h6310d30d;
	16'h1e66 : data <= 32'h13020000;
	16'h1e67 : data <= 32'hb710f00f;
	16'h1e68 : data <= 32'h938000ff;
	16'h1e69 : data <= 32'h93c1000f;
	16'h1e6a : data <= 32'h13021200;
	16'h1e6b : data <= 32'h93022000;
	16'h1e6c : data <= 32'he31652fe;
	16'h1e6d : data <= 32'hb71ef00f;
	16'h1e6e : data <= 32'h938e0ef0;
	16'h1e6f : data <= 32'h130e4030;
	16'h1e70 : data <= 32'h639ad109;
	16'h1e71 : data <= 32'h13020000;
	16'h1e72 : data <= 32'hb710ff00;
	16'h1e73 : data <= 32'h9380f0ff;
	16'h1e74 : data <= 32'h13000000;
	16'h1e75 : data <= 32'h93c1f000;
	16'h1e76 : data <= 32'h13021200;
	16'h1e77 : data <= 32'h93022000;
	16'h1e78 : data <= 32'he31452fe;
	16'h1e79 : data <= 32'hb71eff00;
	16'h1e7a : data <= 32'h938e0eff;
	16'h1e7b : data <= 32'h130e5030;
	16'h1e7c : data <= 32'h6392d107;
	16'h1e7d : data <= 32'h13020000;
	16'h1e7e : data <= 32'hb7f00ff0;
	16'h1e7f : data <= 32'h9380f000;
	16'h1e80 : data <= 32'h13000000;
	16'h1e81 : data <= 32'h13000000;
	16'h1e82 : data <= 32'h93c1000f;
	16'h1e83 : data <= 32'h13021200;
	16'h1e84 : data <= 32'h93022000;
	16'h1e85 : data <= 32'he31252fe;
	16'h1e86 : data <= 32'hb7fe0ff0;
	16'h1e87 : data <= 32'h938efe0f;
	16'h1e88 : data <= 32'h130e6030;
	16'h1e89 : data <= 32'h6398d103;
	16'h1e8a : data <= 32'h9340000f;
	16'h1e8b : data <= 32'h930e000f;
	16'h1e8c : data <= 32'h130e7030;
	16'h1e8d : data <= 32'h6390d003;
	16'h1e8e : data <= 32'hb700ff00;
	16'h1e8f : data <= 32'h9380f00f;
	16'h1e90 : data <= 32'h13c0f070;
	16'h1e91 : data <= 32'h930e0000;
	16'h1e92 : data <= 32'h130e8030;
	16'h1e93 : data <= 32'h6314d001;
	16'h1e94 : data <= 32'h631cc001;
	16'h1e95 : data <= 32'h0f00f00f;
	16'h1e96 : data <= 32'h63000e00;
	16'h1e97 : data <= 32'h131e1e00;
	16'h1e98 : data <= 32'h136e1e00;
	16'h1e99 : data <= 32'h6f000001;
	16'h1e9a : data <= 32'h0f00f00f;
	16'h1e9b : data <= 32'h130e1000;
	16'h1e9c : data <= 32'h6f004000;
	16'h1e9d : data <= 32'h8322c00f;
	16'h1e9e : data <= 32'h1303e003;
	16'h1e9f : data <= 32'hb3035340;
	16'h1ea0 : data <= 32'hb3837300;
	16'h1ea1 : data <= 32'hb3837300;
	16'h1ea2 : data <= 32'h23247000;
	16'h1ea3 : data <= 32'h83228000;
	16'h1ea4 : data <= 32'h13834200;
	16'h1ea5 : data <= 32'h23246000;
	16'h1ea6 : data <= 32'h9303c00f;
	16'h1ea7 : data <= 32'h63147300;
	16'h1ea8 : data <= 32'h6f000000;
	16'h1ea9 : data <= 32'h2322c001;
	16'h1eaa : data <= 32'h83238000;
	16'h1eab : data <= 32'h03a30300;
	16'h1eac : data <= 32'h93034300;
	16'h1ead : data <= 32'h23267000;
	16'h1eae : data <= 32'h67000300;
	16'h1eaf : data <= 32'hff00f00f;
	16'h1eb0 : data <= 32'hff00f00f;
	16'h1eb1 : data <= 32'hff0000ff;
	16'h1eb2 : data <= 32'hf00f0ff0;
	16'h1eb3 : data <= 32'hff0000ff;
	16'h1eb4 : data <= 32'hf00f0ff0;
	16'h1eb5 : data <= 32'hff00ff00;
	16'h1eb6 : data <= 32'h00ff00ff;
	16'h1eb7 : data <= 32'hf00ff00f;
	16'h1eb8 : data <= 32'h0ff00ff0;
	16'h1eb9 : data <= 32'hefefefef;
	16'h1eba : data <= 32'hefefefef;
	16'h1ebb : data <= 32'hefefefbe;
	16'h1ebc : data <= 32'hefbeefbe;
	16'h1ebd : data <= 32'hefbeefbe;
	16'h1ebe : data <= 32'hefbeefbe;
	16'h1ebf : data <= 32'hefbeefbe;
	16'h1ec0 : data <= 32'hefbeefbe;
	16'h1ec1 : data <= 32'haddeefbe;
	16'h1ec2 : data <= 32'haddeefbe;
	16'h1ec3 : data <= 32'haddeefbe;
	16'h1ec4 : data <= 32'haddeefbe;
	16'h1ec5 : data <= 32'haddeefbe;
	16'h1ec6 : data <= 32'haddeefbe;
	16'h1ec7 : data <= 32'haddeefbe;
	16'h1ec8 : data <= 32'haddeefbe;
	16'h1ec9 : data <= 32'haddeefbe;
	16'h1eca : data <= 32'hadde0000;
	16'h1ecb : data <= 32'hFF;
	16'h3c : data <= 32'h307c0000;
	16'h1ecc : data <= 32'h13000000;
	16'h1ecd : data <= 32'h13000000;
	16'h1ece : data <= 32'h13000000;
	16'h1ecf : data <= 32'h13000000;
	16'h1ed0 : data <= 32'h13000000;
	16'h1ed1 : data <= 32'h13000000;
	16'h1ed2 : data <= 32'h13000000;
	16'h1ed3 : data <= 32'h13000000;
	16'h1ed4 : data <= 32'h13000000;
	16'h1ed5 : data <= 32'h13000000;
	16'h1ed6 : data <= 32'h13000000;
	16'h1ed7 : data <= 32'h13000000;
	16'h1ed8 : data <= 32'h13000000;
	16'h1ed9 : data <= 32'h13000000;
	16'h1eda : data <= 32'h13000000;
	16'h1edb : data <= 32'h13000000;
	16'h1edc : data <= 32'h13000000;
	16'h1edd : data <= 32'h13000000;
	16'h1ede : data <= 32'h13000000;
	16'h1edf : data <= 32'h13000000;
	16'h1ee0 : data <= 32'h13000000;
	16'h1ee1 : data <= 32'h13000000;
	16'h1ee2 : data <= 32'h13000000;
	16'h1ee3 : data <= 32'h13000000;
	16'h1ee4 : data <= 32'h13000000;
	16'h1ee5 : data <= 32'h13000000;
	16'h1ee6 : data <= 32'h13000000;
	16'h1ee7 : data <= 32'h13000000;
	16'h1ee8 : data <= 32'h13000000;
	16'h1ee9 : data <= 32'h13000000;
	16'h1eea : data <= 32'h13000000;
	16'h1eeb : data <= 32'h13000000;
	16'h1eec : data <= 32'h13000000;
	16'h1eed : data <= 32'h13000000;
	16'h1eee : data <= 32'h13000000;
	16'h1eef : data <= 32'h13000000;
	16'h1ef0 : data <= 32'h13000000;
	16'h1ef1 : data <= 32'h13000000;
	16'h1ef2 : data <= 32'h13000000;
	16'h1ef3 : data <= 32'h13000000;
	16'h1ef4 : data <= 32'h13000000;
	16'h1ef5 : data <= 32'h13000000;
	16'h1ef6 : data <= 32'h13000000;
	16'h1ef7 : data <= 32'h13000000;
	16'h1ef8 : data <= 32'h13000000;
	16'h1ef9 : data <= 32'h13000000;
	16'h1efa : data <= 32'h13000000;
	16'h1efb : data <= 32'h13000000;
	16'h1efc : data <= 32'h1301c1ff;
	16'h1efd : data <= 32'h23201100;
	16'h1efe : data <= 32'hef004006;
	16'h1eff : data <= 32'h83200100;
	16'h1f00 : data <= 32'h13014100;
	16'h1f01 : data <= 32'h73000010;
	16'h1f02 : data <= 32'h13000000;
	16'h1f03 : data <= 32'h13000000;
	16'h1f04 : data <= 32'h13000000;
	16'h1f05 : data <= 32'h13000000;
	16'h1f06 : data <= 32'h13000000;
	16'h1f07 : data <= 32'h13000000;
	16'h1f08 : data <= 32'h13000000;
	16'h1f09 : data <= 32'h13000000;
	16'h1f0a : data <= 32'h13000000;
	16'h1f0b : data <= 32'h13000000;
	16'h1f0c : data <= 32'h13610000;
	16'h1f0d : data <= 32'h1301c1ff;
	16'h1f0e : data <= 32'h9362c000;
	16'h1f0f : data <= 32'h9392c201;
	16'h1f10 : data <= 32'h13630000;
	16'h1f11 : data <= 32'h1303f3ff;
	16'h1f12 : data <= 32'hb3c26200;
	16'h1f13 : data <= 32'h33715100;
	16'h1f14 : data <= 32'h97020000;
	16'h1f15 : data <= 32'h9382c27a;
	16'h1f16 : data <= 32'h67800200;
	16'h1f17 : data <= 32'h1301c1ff;
	16'h1f18 : data <= 32'h23201100;
	16'h1f19 : data <= 32'h232ef1ff;
	16'h1f1a : data <= 32'h232ce1ff;
	16'h1f1b : data <= 32'h232ad1ff;
	16'h1f1c : data <= 32'h2328c1ff;
	16'h1f1d : data <= 32'h2326b1ff;
	16'h1f1e : data <= 32'h2324a1ff;
	16'h1f1f : data <= 32'h232291ff;
	16'h1f20 : data <= 32'h232081ff;
	16'h1f21 : data <= 32'h232e71fd;
	16'h1f22 : data <= 32'h232c61fd;
	16'h1f23 : data <= 32'h232a51fd;
	16'h1f24 : data <= 32'h232841fd;
	16'h1f25 : data <= 32'h232631fd;
	16'h1f26 : data <= 32'h232421fd;
	16'h1f27 : data <= 32'h232211fd;
	16'h1f28 : data <= 32'h232001fd;
	16'h1f29 : data <= 32'h232ef1fa;
	16'h1f2a : data <= 32'h232ce1fa;
	16'h1f2b : data <= 32'h232ad1fa;
	16'h1f2c : data <= 32'h2328c1fa;
	16'h1f2d : data <= 32'h2326b1fa;
	16'h1f2e : data <= 32'h2324a1fa;
	16'h1f2f : data <= 32'h232291fa;
	16'h1f30 : data <= 32'h232081fa;
	16'h1f31 : data <= 32'h232e71f8;
	16'h1f32 : data <= 32'h232c61f8;
	16'h1f33 : data <= 32'h232a51f8;
	16'h1f34 : data <= 32'h232841f8;
	16'h1f35 : data <= 32'h232631f8;
	16'h1f36 : data <= 32'h232421f8;
	16'h1f37 : data <= 32'h232211f8;
	16'h1f38 : data <= 32'h232001f8;
	16'h1f39 : data <= 32'h130101f8;
	16'h1f3a : data <= 32'h93050100;
	16'h1f3b : data <= 32'h73261034;
	16'h1f3c : data <= 32'hf3263034;
	16'h1f3d : data <= 32'h73252034;
	16'h1f3e : data <= 32'h93020500;
	16'h1f3f : data <= 32'h93d2f201;
	16'h1f40 : data <= 32'h63860200;
	16'h1f41 : data <= 32'hef004009;
	16'h1f42 : data <= 32'h6f004001;
	16'h1f43 : data <= 32'hef00400d;
	16'h1f44 : data <= 32'hf3221034;
	16'h1f45 : data <= 32'h93824200;
	16'h1f46 : data <= 32'h73901234;
	16'h1f47 : data <= 32'h832fc107;
	16'h1f48 : data <= 32'h032f8107;
	16'h1f49 : data <= 32'h832e4107;
	16'h1f4a : data <= 32'h032e0107;
	16'h1f4b : data <= 32'h832dc106;
	16'h1f4c : data <= 32'h032d8106;
	16'h1f4d : data <= 32'h832c4106;
	16'h1f4e : data <= 32'h032c0106;
	16'h1f4f : data <= 32'h832bc105;
	16'h1f50 : data <= 32'h032b8105;
	16'h1f51 : data <= 32'h832a4105;
	16'h1f52 : data <= 32'h032a0105;
	16'h1f53 : data <= 32'h8329c104;
	16'h1f54 : data <= 32'h03298104;
	16'h1f55 : data <= 32'h83284104;
	16'h1f56 : data <= 32'h03280104;
	16'h1f57 : data <= 32'h8327c103;
	16'h1f58 : data <= 32'h03278103;
	16'h1f59 : data <= 32'h83264103;
	16'h1f5a : data <= 32'h03260103;
	16'h1f5b : data <= 32'h8325c102;
	16'h1f5c : data <= 32'h03258102;
	16'h1f5d : data <= 32'h83244102;
	16'h1f5e : data <= 32'h03240102;
	16'h1f5f : data <= 32'h8323c101;
	16'h1f60 : data <= 32'h03238101;
	16'h1f61 : data <= 32'h83224101;
	16'h1f62 : data <= 32'h13010108;
	16'h1f63 : data <= 32'h83200100;
	16'h1f64 : data <= 32'h13014100;
	16'h1f65 : data <= 32'h67800000;
	16'h1f66 : data <= 32'h130101fe;
	16'h1f67 : data <= 32'h232e8100;
	16'h1f68 : data <= 32'h13040102;
	16'h1f69 : data <= 32'h2326a4fe;
	16'h1f6a : data <= 32'h13000000;
	16'h1f6b : data <= 32'h0324c101;
	16'h1f6c : data <= 32'h13010102;
	16'h1f6d : data <= 32'h67800000;
	16'h1f6e : data <= 32'h130101fe;
	16'h1f6f : data <= 32'h232e8100;
	16'h1f70 : data <= 32'h13040102;
	16'h1f71 : data <= 32'h2326a4fe;
	16'h1f72 : data <= 32'h8327c4fe;
	16'h1f73 : data <= 32'hb307f040;
	16'h1f74 : data <= 32'h13850700;
	16'h1f75 : data <= 32'h0324c101;
	16'h1f76 : data <= 32'h13010102;
	16'h1f77 : data <= 32'h67800000;
	16'h1f78 : data <= 32'h130101fb;
	16'h1f79 : data <= 32'h23261104;
	16'h1f7a : data <= 32'h23248104;
	16'h1f7b : data <= 32'h23229104;
	16'h1f7c : data <= 32'h13040105;
	16'h1f7d : data <= 32'h232ea4fa;
	16'h1f7e : data <= 32'h232cb4fa;
	16'h1f7f : data <= 32'h232ac4fa;
	16'h1f80 : data <= 32'h2328d4fa;
	16'h1f81 : data <= 32'h0327c4fb;
	16'h1f82 : data <= 32'h93072000;
	16'h1f83 : data <= 32'h6312f752;
	16'h1f84 : data <= 32'h832744fb;
	16'h1f85 : data <= 32'h83a70700;
	16'h1f86 : data <= 32'h2326f4fe;
	16'h1f87 : data <= 32'h8327c4fe;
	16'h1f88 : data <= 32'h93f7f707;
	16'h1f89 : data <= 32'h2324f4fe;
	16'h1f8a : data <= 32'h0327c4fe;
	16'h1f8b : data <= 32'hb7170000;
	16'h1f8c : data <= 32'h938707f8;
	16'h1f8d : data <= 32'hb377f700;
	16'h1f8e : data <= 32'h93d77740;
	16'h1f8f : data <= 32'h2322f4fe;
	16'h1f90 : data <= 32'h0327c4fe;
	16'h1f91 : data <= 32'hb7870f00;
	16'h1f92 : data <= 32'hb377f700;
	16'h1f93 : data <= 32'h93d7f740;
	16'h1f94 : data <= 32'h2320f4fe;
	16'h1f95 : data <= 32'h0327c4fe;
	16'h1f96 : data <= 32'hb707f001;
	16'h1f97 : data <= 32'hb377f700;
	16'h1f98 : data <= 32'h93d74741;
	16'h1f99 : data <= 32'h232ef4fc;
	16'h1f9a : data <= 32'h0327c4fe;
	16'h1f9b : data <= 32'hb7770000;
	16'h1f9c : data <= 32'hb377f700;
	16'h1f9d : data <= 32'h93d7c740;
	16'h1f9e : data <= 32'h232cf4fc;
	16'h1f9f : data <= 32'h8327c4fe;
	16'h1fa0 : data <= 32'h93d79701;
	16'h1fa1 : data <= 32'h232af4fc;
	16'h1fa2 : data <= 32'h032784fe;
	16'h1fa3 : data <= 32'h93073003;
	16'h1fa4 : data <= 32'h6310f74a;
	16'h1fa5 : data <= 32'h032744fd;
	16'h1fa6 : data <= 32'h93071000;
	16'h1fa7 : data <= 32'h631af748;
	16'h1fa8 : data <= 32'h832784fd;
	16'h1fa9 : data <= 32'h63960704;
	16'h1faa : data <= 32'h8327c4fd;
	16'h1fab : data <= 32'h93972700;
	16'h1fac : data <= 32'h032784fb;
	16'h1fad : data <= 32'hb307f700;
	16'h1fae : data <= 32'h83a60700;
	16'h1faf : data <= 32'h832704fe;
	16'h1fb0 : data <= 32'h93972700;
	16'h1fb1 : data <= 32'h032784fb;
	16'h1fb2 : data <= 32'hb307f700;
	16'h1fb3 : data <= 32'h83a50700;
	16'h1fb4 : data <= 32'h832744fe;
	16'h1fb5 : data <= 32'h93972700;
	16'h1fb6 : data <= 32'h032784fb;
	16'h1fb7 : data <= 32'hb307f700;
	16'h1fb8 : data <= 32'h13860700;
	16'h1fb9 : data <= 32'h13850600;
	16'h1fba : data <= 32'hef000046;
	16'h1fbb : data <= 32'h6f004044;
	16'h1fbc : data <= 32'h032784fd;
	16'h1fbd : data <= 32'h93071000;
	16'h1fbe : data <= 32'h630cf742;
	16'h1fbf : data <= 32'h032784fd;
	16'h1fc0 : data <= 32'h93072000;
	16'h1fc1 : data <= 32'h6306f742;
	16'h1fc2 : data <= 32'h032784fd;
	16'h1fc3 : data <= 32'h93073000;
	16'h1fc4 : data <= 32'h6300f742;
	16'h1fc5 : data <= 32'h032784fd;
	16'h1fc6 : data <= 32'h93074000;
	16'h1fc7 : data <= 32'h631cf716;
	16'h1fc8 : data <= 32'h8327c4fd;
	16'h1fc9 : data <= 32'h93972700;
	16'h1fca : data <= 32'h032784fb;
	16'h1fcb : data <= 32'hb307f700;
	16'h1fcc : data <= 32'h83a70700;
	16'h1fcd : data <= 32'h2328f4fc;
	16'h1fce : data <= 32'h832704fe;
	16'h1fcf : data <= 32'h93972700;
	16'h1fd0 : data <= 32'h032784fb;
	16'h1fd1 : data <= 32'hb307f700;
	16'h1fd2 : data <= 32'h83a70700;
	16'h1fd3 : data <= 32'h2326f4fc;
	16'h1fd4 : data <= 32'h832704fd;
	16'h1fd5 : data <= 32'h639c0700;
	16'h1fd6 : data <= 32'h9307f0ff;
	16'h1fd7 : data <= 32'h2324f4fc;
	16'h1fd8 : data <= 32'h8327c4fc;
	16'h1fd9 : data <= 32'h2322f4fc;
	16'h1fda : data <= 32'h6f000011;
	16'h1fdb : data <= 32'h0327c4fc;
	16'h1fdc : data <= 32'hb7070080;
	16'h1fdd : data <= 32'h6310f702;
	16'h1fde : data <= 32'h032704fd;
	16'h1fdf : data <= 32'h9307f0ff;
	16'h1fe0 : data <= 32'h631af700;
	16'h1fe1 : data <= 32'h8327c4fc;
	16'h1fe2 : data <= 32'h2324f4fc;
	16'h1fe3 : data <= 32'h232204fc;
	16'h1fe4 : data <= 32'h6f00800e;
	16'h1fe5 : data <= 32'h8327c4fc;
	16'h1fe6 : data <= 32'h63d00704;
	16'h1fe7 : data <= 32'h832704fd;
	16'h1fe8 : data <= 32'h63dc0702;
	16'h1fe9 : data <= 32'h0325c4fc;
	16'h1fea : data <= 32'heff01fe1;
	16'h1feb : data <= 32'h93040500;
	16'h1fec : data <= 32'h032504fd;
	16'h1fed : data <= 32'heff05fe0;
	16'h1fee : data <= 32'h93050500;
	16'h1fef : data <= 32'h130744fc;
	16'h1ff0 : data <= 32'h930784fc;
	16'h1ff1 : data <= 32'h93060700;
	16'h1ff2 : data <= 32'h13860700;
	16'h1ff3 : data <= 32'h13850400;
	16'h1ff4 : data <= 32'hef00403c;
	16'h1ff5 : data <= 32'h6f00400a;
	16'h1ff6 : data <= 32'h8327c4fc;
	16'h1ff7 : data <= 32'h63de0702;
	16'h1ff8 : data <= 32'h0325c4fc;
	16'h1ff9 : data <= 32'heff05fdd;
	16'h1ffa : data <= 32'h130744fc;
	16'h1ffb : data <= 32'h930784fc;
	16'h1ffc : data <= 32'h93060700;
	16'h1ffd : data <= 32'h13860700;
	16'h1ffe : data <= 32'h832504fd;
	16'h1fff : data <= 32'hef008039;
	16'h2000 : data <= 32'h832784fc;
	16'h2001 : data <= 32'h13850700;
	16'h2002 : data <= 32'heff01fdb;
	16'h2003 : data <= 32'h93070500;
	16'h2004 : data <= 32'h2324f4fc;
	16'h2005 : data <= 32'h6f004006;
	16'h2006 : data <= 32'h832704fd;
	16'h2007 : data <= 32'h63d00704;
	16'h2008 : data <= 32'h032504fd;
	16'h2009 : data <= 32'heff05fd9;
	16'h200a : data <= 32'h93050500;
	16'h200b : data <= 32'h130744fc;
	16'h200c : data <= 32'h930784fc;
	16'h200d : data <= 32'h93060700;
	16'h200e : data <= 32'h13860700;
	16'h200f : data <= 32'h0325c4fc;
	16'h2010 : data <= 32'hef004035;
	16'h2011 : data <= 32'h832784fc;
	16'h2012 : data <= 32'h13850700;
	16'h2013 : data <= 32'heff0dfd6;
	16'h2014 : data <= 32'h93070500;
	16'h2015 : data <= 32'h2324f4fc;
	16'h2016 : data <= 32'h6f000002;
	16'h2017 : data <= 32'h130744fc;
	16'h2018 : data <= 32'h930784fc;
	16'h2019 : data <= 32'h93060700;
	16'h201a : data <= 32'h13860700;
	16'h201b : data <= 32'h832504fd;
	16'h201c : data <= 32'h0325c4fc;
	16'h201d : data <= 32'hef000032;
	16'h201e : data <= 32'h832744fe;
	16'h201f : data <= 32'h93972700;
	16'h2020 : data <= 32'h032784fb;
	16'h2021 : data <= 32'hb307f700;
	16'h2022 : data <= 32'h032784fc;
	16'h2023 : data <= 32'h23a0e700;
	16'h2024 : data <= 32'h6f00002a;
	16'h2025 : data <= 32'h032784fd;
	16'h2026 : data <= 32'h93075000;
	16'h2027 : data <= 32'h6314f708;
	16'h2028 : data <= 32'h8327c4fd;
	16'h2029 : data <= 32'h93972700;
	16'h202a : data <= 32'h032784fb;
	16'h202b : data <= 32'hb307f700;
	16'h202c : data <= 32'h83a70700;
	16'h202d : data <= 32'h2328f4fc;
	16'h202e : data <= 32'h832704fe;
	16'h202f : data <= 32'h93972700;
	16'h2030 : data <= 32'h032784fb;
	16'h2031 : data <= 32'hb307f700;
	16'h2032 : data <= 32'h83a70700;
	16'h2033 : data <= 32'h2326f4fc;
	16'h2034 : data <= 32'h832704fd;
	16'h2035 : data <= 32'h639c0700;
	16'h2036 : data <= 32'h9307f0ff;
	16'h2037 : data <= 32'h2324f4fc;
	16'h2038 : data <= 32'h8327c4fc;
	16'h2039 : data <= 32'h2322f4fc;
	16'h203a : data <= 32'h6f000002;
	16'h203b : data <= 32'h130744fc;
	16'h203c : data <= 32'h930784fc;
	16'h203d : data <= 32'h93060700;
	16'h203e : data <= 32'h13860700;
	16'h203f : data <= 32'h832504fd;
	16'h2040 : data <= 32'h0325c4fc;
	16'h2041 : data <= 32'hef000029;
	16'h2042 : data <= 32'h832744fe;
	16'h2043 : data <= 32'h93972700;
	16'h2044 : data <= 32'h032784fb;
	16'h2045 : data <= 32'hb307f700;
	16'h2046 : data <= 32'h032784fc;
	16'h2047 : data <= 32'h23a0e700;
	16'h2048 : data <= 32'h6f000021;
	16'h2049 : data <= 32'h032784fd;
	16'h204a : data <= 32'h93076000;
	16'h204b : data <= 32'h631cf716;
	16'h204c : data <= 32'h8327c4fd;
	16'h204d : data <= 32'h93972700;
	16'h204e : data <= 32'h032784fb;
	16'h204f : data <= 32'hb307f700;
	16'h2050 : data <= 32'h83a70700;
	16'h2051 : data <= 32'h2328f4fc;
	16'h2052 : data <= 32'h832704fe;
	16'h2053 : data <= 32'h93972700;
	16'h2054 : data <= 32'h032784fb;
	16'h2055 : data <= 32'hb307f700;
	16'h2056 : data <= 32'h83a70700;
	16'h2057 : data <= 32'h2326f4fc;
	16'h2058 : data <= 32'h832704fd;
	16'h2059 : data <= 32'h639c0700;
	16'h205a : data <= 32'h9307f0ff;
	16'h205b : data <= 32'h2324f4fc;
	16'h205c : data <= 32'h8327c4fc;
	16'h205d : data <= 32'h2322f4fc;
	16'h205e : data <= 32'h6f000011;
	16'h205f : data <= 32'h0327c4fc;
	16'h2060 : data <= 32'hb7070080;
	16'h2061 : data <= 32'h6310f702;
	16'h2062 : data <= 32'h032704fd;
	16'h2063 : data <= 32'h9307f0ff;
	16'h2064 : data <= 32'h631af700;
	16'h2065 : data <= 32'h8327c4fc;
	16'h2066 : data <= 32'h2324f4fc;
	16'h2067 : data <= 32'h232204fc;
	16'h2068 : data <= 32'h6f00800e;
	16'h2069 : data <= 32'h8327c4fc;
	16'h206a : data <= 32'h63d00704;
	16'h206b : data <= 32'h832704fd;
	16'h206c : data <= 32'h63dc0702;
	16'h206d : data <= 32'h0325c4fc;
	16'h206e : data <= 32'heff01fc0;
	16'h206f : data <= 32'h93040500;
	16'h2070 : data <= 32'h032504fd;
	16'h2071 : data <= 32'heff05fbf;
	16'h2072 : data <= 32'h93050500;
	16'h2073 : data <= 32'h130744fc;
	16'h2074 : data <= 32'h930784fc;
	16'h2075 : data <= 32'h93060700;
	16'h2076 : data <= 32'h13860700;
	16'h2077 : data <= 32'h13850400;
	16'h2078 : data <= 32'hef00401b;
	16'h2079 : data <= 32'h6f00400a;
	16'h207a : data <= 32'h8327c4fc;
	16'h207b : data <= 32'h63de0702;
	16'h207c : data <= 32'h0325c4fc;
	16'h207d : data <= 32'heff05fbc;
	16'h207e : data <= 32'h130744fc;
	16'h207f : data <= 32'h930784fc;
	16'h2080 : data <= 32'h93060700;
	16'h2081 : data <= 32'h13860700;
	16'h2082 : data <= 32'h832504fd;
	16'h2083 : data <= 32'hef008018;
	16'h2084 : data <= 32'h832744fc;
	16'h2085 : data <= 32'h13850700;
	16'h2086 : data <= 32'heff01fba;
	16'h2087 : data <= 32'h93070500;
	16'h2088 : data <= 32'h2322f4fc;
	16'h2089 : data <= 32'h6f004006;
	16'h208a : data <= 32'h832704fd;
	16'h208b : data <= 32'h63d00704;
	16'h208c : data <= 32'h032504fd;
	16'h208d : data <= 32'heff05fb8;
	16'h208e : data <= 32'h93050500;
	16'h208f : data <= 32'h130744fc;
	16'h2090 : data <= 32'h930784fc;
	16'h2091 : data <= 32'h93060700;
	16'h2092 : data <= 32'h13860700;
	16'h2093 : data <= 32'h0325c4fc;
	16'h2094 : data <= 32'hef004014;
	16'h2095 : data <= 32'h832744fc;
	16'h2096 : data <= 32'h13850700;
	16'h2097 : data <= 32'heff0dfb5;
	16'h2098 : data <= 32'h93070500;
	16'h2099 : data <= 32'h2322f4fc;
	16'h209a : data <= 32'h6f000002;
	16'h209b : data <= 32'h130744fc;
	16'h209c : data <= 32'h930784fc;
	16'h209d : data <= 32'h93060700;
	16'h209e : data <= 32'h13860700;
	16'h209f : data <= 32'h832504fd;
	16'h20a0 : data <= 32'h0325c4fc;
	16'h20a1 : data <= 32'hef000011;
	16'h20a2 : data <= 32'h832744fe;
	16'h20a3 : data <= 32'h93972700;
	16'h20a4 : data <= 32'h032784fb;
	16'h20a5 : data <= 32'hb307f700;
	16'h20a6 : data <= 32'h032744fc;
	16'h20a7 : data <= 32'h23a0e700;
	16'h20a8 : data <= 32'h6f000009;
	16'h20a9 : data <= 32'h032784fd;
	16'h20aa : data <= 32'h93077000;
	16'h20ab : data <= 32'h6312f708;
	16'h20ac : data <= 32'h8327c4fd;
	16'h20ad : data <= 32'h93972700;
	16'h20ae : data <= 32'h032784fb;
	16'h20af : data <= 32'hb307f700;
	16'h20b0 : data <= 32'h83a70700;
	16'h20b1 : data <= 32'h2328f4fc;
	16'h20b2 : data <= 32'h832704fe;
	16'h20b3 : data <= 32'h93972700;
	16'h20b4 : data <= 32'h032784fb;
	16'h20b5 : data <= 32'hb307f700;
	16'h20b6 : data <= 32'h83a70700;
	16'h20b7 : data <= 32'h2326f4fc;
	16'h20b8 : data <= 32'h832704fd;
	16'h20b9 : data <= 32'h639c0700;
	16'h20ba : data <= 32'h9307f0ff;
	16'h20bb : data <= 32'h2324f4fc;
	16'h20bc : data <= 32'h8327c4fc;
	16'h20bd : data <= 32'h2322f4fc;
	16'h20be : data <= 32'h6f000002;
	16'h20bf : data <= 32'h130744fc;
	16'h20c0 : data <= 32'h930784fc;
	16'h20c1 : data <= 32'h93060700;
	16'h20c2 : data <= 32'h13860700;
	16'h20c3 : data <= 32'h832504fd;
	16'h20c4 : data <= 32'h0325c4fc;
	16'h20c5 : data <= 32'hef000008;
	16'h20c6 : data <= 32'h832744fe;
	16'h20c7 : data <= 32'h93972700;
	16'h20c8 : data <= 32'h032784fb;
	16'h20c9 : data <= 32'hb307f700;
	16'h20ca : data <= 32'h032744fc;
	16'h20cb : data <= 32'h23a0e700;
	16'h20cc : data <= 32'h13000000;
	16'h20cd : data <= 32'h8320c104;
	16'h20ce : data <= 32'h03248104;
	16'h20cf : data <= 32'h83244104;
	16'h20d0 : data <= 32'h13010105;
	16'h20d1 : data <= 32'h67800000;
	16'h20d2 : data <= 32'h130101fe;
	16'h20d3 : data <= 32'h232e8100;
	16'h20d4 : data <= 32'h13040102;
	16'h20d5 : data <= 32'h2326a4fe;
	16'h20d6 : data <= 32'h2324b4fe;
	16'h20d7 : data <= 32'h2322c4fe;
	16'h20d8 : data <= 32'h93020500;
	16'h20d9 : data <= 32'h13050000;
	16'h20da : data <= 32'h13f31500;
	16'h20db : data <= 32'h63040300;
	16'h20dc : data <= 32'h3385a200;
	16'h20dd : data <= 32'h93921200;
	16'h20de : data <= 32'h93d51500;
	16'h20df : data <= 32'he39605fe;
	16'h20e0 : data <= 32'h2320a600;
	16'h20e1 : data <= 32'h13000000;
	16'h20e2 : data <= 32'h0324c101;
	16'h20e3 : data <= 32'h13010102;
	16'h20e4 : data <= 32'h67800000;
	16'h20e5 : data <= 32'h130101fe;
	16'h20e6 : data <= 32'h232e8100;
	16'h20e7 : data <= 32'h13040102;
	16'h20e8 : data <= 32'h2326a4fe;
	16'h20e9 : data <= 32'h2324b4fe;
	16'h20ea : data <= 32'h2322c4fe;
	16'h20eb : data <= 32'h2320d4fe;
	16'h20ec : data <= 32'h93020000;
	16'h20ed : data <= 32'h13030000;
	16'h20ee : data <= 32'h130e1000;
	16'h20ef : data <= 32'h131efe01;
	16'h20f0 : data <= 32'h13131300;
	16'h20f1 : data <= 32'hb373c501;
	16'h20f2 : data <= 32'h63840300;
	16'h20f3 : data <= 32'h13631300;
	16'h20f4 : data <= 32'h6346b300;
	16'h20f5 : data <= 32'h3303b340;
	16'h20f6 : data <= 32'hb3e2c201;
	16'h20f7 : data <= 32'h135e1e00;
	16'h20f8 : data <= 32'he3100efe;
	16'h20f9 : data <= 32'h23205600;
	16'h20fa : data <= 32'h23a06600;
	16'h20fb : data <= 32'h13000000;
	16'h20fc : data <= 32'h0324c101;
	16'h20fd : data <= 32'h13010102;
	16'h20fe : data <= 32'h67800000;
	16'h20ff : data <= 32'h130101ff;
	16'h2100 : data <= 32'h23268100;
	16'h2101 : data <= 32'h13040101;
	16'h2102 : data <= 32'h83228000;
	16'h2103 : data <= 32'h13834200;
	16'h2104 : data <= 32'h23246000;
	16'h2105 : data <= 32'h9303c00f;
	16'h2106 : data <= 32'h63147300;
	16'h2107 : data <= 32'h6f000000;
	16'h2108 : data <= 32'h83238000;
	16'h2109 : data <= 32'h03a30300;
	16'h210a : data <= 32'h67000300;
	16'h210b : data <= 32'h13000000;
	16'h210c : data <= 32'h13850700;
	16'h210d : data <= 32'h0324c100;
	16'h210e : data <= 32'h13010101;
	16'h210f : data <= 32'h67800000;
	16'h2110 : data <= 32'h130101fd;
	16'h2111 : data <= 32'h23268102;
	16'h2112 : data <= 32'h13040103;
	16'h2113 : data <= 32'h232ea4fc;
	16'h2114 : data <= 32'h232cb4fc;
	16'h2115 : data <= 32'h232ac4fc;
	16'h2116 : data <= 32'h2328d4fc;
	16'h2117 : data <= 32'h8327c4fd;
	16'h2118 : data <= 32'h83a70700;
	16'h2119 : data <= 32'h032784fd;
	16'h211a : data <= 32'h23a4e700;
	16'h211b : data <= 32'h8327c4fd;
	16'h211c : data <= 32'h83a70700;
	16'h211d : data <= 32'h032704fd;
	16'h211e : data <= 32'h23aae700;
	16'h211f : data <= 32'h8327c4fd;
	16'h2120 : data <= 32'h83a70700;
	16'h2121 : data <= 32'h83a74700;
	16'h2122 : data <= 32'h2326f4fe;
	16'h2123 : data <= 32'h8327c4fe;
	16'h2124 : data <= 32'h93f7e7ff;
	16'h2125 : data <= 32'h2326f4fe;
	16'h2126 : data <= 32'h8327c4fd;
	16'h2127 : data <= 32'h83a70700;
	16'h2128 : data <= 32'h032744fd;
	16'h2129 : data <= 32'h93761700;
	16'h212a : data <= 32'h0327c4fe;
	16'h212b : data <= 32'h33e7e600;
	16'h212c : data <= 32'h23a2e700;
	16'h212d : data <= 32'h93070000;
	16'h212e : data <= 32'h13850700;
	16'h212f : data <= 32'h0324c102;
	16'h2130 : data <= 32'h13010103;
	16'h2131 : data <= 32'h67800000;
	16'h2132 : data <= 32'h130101fc;
	16'h2133 : data <= 32'h232e8102;
	16'h2134 : data <= 32'h13040104;
	16'h2135 : data <= 32'h2326a4fc;
	16'h2136 : data <= 32'h2324b4fc;
	16'h2137 : data <= 32'h2322c4fc;
	16'h2138 : data <= 32'h232604fe;
	16'h2139 : data <= 32'h032744fc;
	16'h213a : data <= 32'h93070004;
	16'h213b : data <= 32'h63f6e700;
	16'h213c : data <= 32'h93070003;
	16'h213d : data <= 32'h6f004020;
	16'h213e : data <= 32'h032744fc;
	16'h213f : data <= 32'h93070004;
	16'h2140 : data <= 32'h631af702;
	16'h2141 : data <= 32'h8327c4fc;
	16'h2142 : data <= 32'h83a70700;
	16'h2143 : data <= 32'h83a74700;
	16'h2144 : data <= 32'h2322f4fe;
	16'h2145 : data <= 32'h832744fe;
	16'h2146 : data <= 32'h93f707fc;
	16'h2147 : data <= 32'h2322f4fe;
	16'h2148 : data <= 32'h8327c4fc;
	16'h2149 : data <= 32'h83a70700;
	16'h214a : data <= 32'h032744fe;
	16'h214b : data <= 32'h23a2e700;
	16'h214c : data <= 32'h6f000004;
	16'h214d : data <= 32'h8327c4fc;
	16'h214e : data <= 32'h83a70700;
	16'h214f : data <= 32'h83a74700;
	16'h2150 : data <= 32'h2320f4fe;
	16'h2151 : data <= 32'h832704fe;
	16'h2152 : data <= 32'h93f707fc;
	16'h2153 : data <= 32'h2320f4fe;
	16'h2154 : data <= 32'h8327c4fc;
	16'h2155 : data <= 32'h83a70700;
	16'h2156 : data <= 32'h032744fc;
	16'h2157 : data <= 32'h13172700;
	16'h2158 : data <= 32'h9376f70f;
	16'h2159 : data <= 32'h032704fe;
	16'h215a : data <= 32'h33e7e600;
	16'h215b : data <= 32'h23a2e700;
	16'h215c : data <= 32'h8327c4fc;
	16'h215d : data <= 32'h83a70700;
	16'h215e : data <= 32'h83a74700;
	16'h215f : data <= 32'h232ef4fc;
	16'h2160 : data <= 32'h8327c4fd;
	16'h2161 : data <= 32'h93f7e7ff;
	16'h2162 : data <= 32'h232ef4fc;
	16'h2163 : data <= 32'h8327c4fc;
	16'h2164 : data <= 32'h83a70700;
	16'h2165 : data <= 32'h0327c4fd;
	16'h2166 : data <= 32'h13670710;
	16'h2167 : data <= 32'h23a2e700;
	16'h2168 : data <= 32'h8327c4fc;
	16'h2169 : data <= 32'h83a70700;
	16'h216a : data <= 32'h83a74700;
	16'h216b : data <= 32'h232cf4fc;
	16'h216c : data <= 32'h832784fd;
	16'h216d : data <= 32'h93f7e7ff;
	16'h216e : data <= 32'h232cf4fc;
	16'h216f : data <= 32'h8327c4fc;
	16'h2170 : data <= 32'h83a70700;
	16'h2171 : data <= 32'h032784fd;
	16'h2172 : data <= 32'h23a2e700;
	16'h2173 : data <= 32'h6f008002;
	16'h2174 : data <= 32'h8327c4fc;
	16'h2175 : data <= 32'h03a70700;
	16'h2176 : data <= 32'h8327c4fe;
	16'h2177 : data <= 32'h93861700;
	16'h2178 : data <= 32'h2326d4fe;
	16'h2179 : data <= 32'h832684fc;
	16'h217a : data <= 32'hb387f600;
	16'h217b : data <= 32'h83c70700;
	16'h217c : data <= 32'h2320f700;
	16'h217d : data <= 32'h0327c4fe;
	16'h217e : data <= 32'h832744fc;
	16'h217f : data <= 32'h637ef700;
	16'h2180 : data <= 32'h8327c4fc;
	16'h2181 : data <= 32'h83a70700;
	16'h2182 : data <= 32'h83a70701;
	16'h2183 : data <= 32'h93d7b700;
	16'h2184 : data <= 32'h93f71700;
	16'h2185 : data <= 32'he38e07fa;
	16'h2186 : data <= 32'h8327c4fc;
	16'h2187 : data <= 32'h83a70700;
	16'h2188 : data <= 32'h83a74700;
	16'h2189 : data <= 32'h232af4fc;
	16'h218a : data <= 32'h832744fd;
	16'h218b : data <= 32'h93f7e7ff;
	16'h218c : data <= 32'h232af4fc;
	16'h218d : data <= 32'h8327c4fc;
	16'h218e : data <= 32'h83a70700;
	16'h218f : data <= 32'h032744fd;
	16'h2190 : data <= 32'h13670720;
	16'h2191 : data <= 32'h23a2e700;
	16'h2192 : data <= 32'h8327c4fc;
	16'h2193 : data <= 32'h83a70700;
	16'h2194 : data <= 32'h83a70701;
	16'h2195 : data <= 32'h2324f4fe;
	16'h2196 : data <= 32'h6f000008;
	16'h2197 : data <= 32'h832784fe;
	16'h2198 : data <= 32'h93f71700;
	16'h2199 : data <= 32'h63860700;
	16'h219a : data <= 32'h93071003;
	16'h219b : data <= 32'h6f00c008;
	16'h219c : data <= 32'h832784fe;
	16'h219d : data <= 32'h93d73700;
	16'h219e : data <= 32'h93f71700;
	16'h219f : data <= 32'h63860700;
	16'h21a0 : data <= 32'h93072003;
	16'h21a1 : data <= 32'h6f004007;
	16'h21a2 : data <= 32'h832784fe;
	16'h21a3 : data <= 32'h93d7b700;
	16'h21a4 : data <= 32'h93f71700;
	16'h21a5 : data <= 32'h639a0702;
	16'h21a6 : data <= 32'h0327c4fe;
	16'h21a7 : data <= 32'h832744fc;
	16'h21a8 : data <= 32'h6374f702;
	16'h21a9 : data <= 32'h8327c4fc;
	16'h21aa : data <= 32'h03a70700;
	16'h21ab : data <= 32'h8327c4fe;
	16'h21ac : data <= 32'h93861700;
	16'h21ad : data <= 32'h2326d4fe;
	16'h21ae : data <= 32'h832684fc;
	16'h21af : data <= 32'hb387f600;
	16'h21b0 : data <= 32'h83c70700;
	16'h21b1 : data <= 32'h2320f700;
	16'h21b2 : data <= 32'h8327c4fc;
	16'h21b3 : data <= 32'h83a70700;
	16'h21b4 : data <= 32'h83a70701;
	16'h21b5 : data <= 32'h2324f4fe;
	16'h21b6 : data <= 32'h0327c4fe;
	16'h21b7 : data <= 32'h832744fc;
	16'h21b8 : data <= 32'he36ef7f6;
	16'h21b9 : data <= 32'h832784fe;
	16'h21ba : data <= 32'h93d72700;
	16'h21bb : data <= 32'h93f71700;
	16'h21bc : data <= 32'he38607f6;
	16'h21bd : data <= 32'h93070000;
	16'h21be : data <= 32'h13850700;
	16'h21bf : data <= 32'h0324c103;
	16'h21c0 : data <= 32'h13010104;
	16'h21c1 : data <= 32'h67800000;
	16'h21c2 : data <= 32'h130101fc;
	16'h21c3 : data <= 32'h232e8102;
	16'h21c4 : data <= 32'h13040104;
	16'h21c5 : data <= 32'h2326a4fc;
	16'h21c6 : data <= 32'h2324b4fc;
	16'h21c7 : data <= 32'h2322c4fc;
	16'h21c8 : data <= 32'h232604fe;
	16'h21c9 : data <= 32'h032744fc;
	16'h21ca : data <= 32'h93070004;
	16'h21cb : data <= 32'h63f6e700;
	16'h21cc : data <= 32'h93070003;
	16'h21cd : data <= 32'h6f00401e;
	16'h21ce : data <= 32'h032744fc;
	16'h21cf : data <= 32'h93070004;
	16'h21d0 : data <= 32'h631af702;
	16'h21d1 : data <= 32'h8327c4fc;
	16'h21d2 : data <= 32'h83a70700;
	16'h21d3 : data <= 32'h83a74700;
	16'h21d4 : data <= 32'h2322f4fe;
	16'h21d5 : data <= 32'h832744fe;
	16'h21d6 : data <= 32'h93f707fc;
	16'h21d7 : data <= 32'h2322f4fe;
	16'h21d8 : data <= 32'h8327c4fc;
	16'h21d9 : data <= 32'h83a70700;
	16'h21da : data <= 32'h032744fe;
	16'h21db : data <= 32'h23a2e700;
	16'h21dc : data <= 32'h6f000004;
	16'h21dd : data <= 32'h8327c4fc;
	16'h21de : data <= 32'h83a70700;
	16'h21df : data <= 32'h83a74700;
	16'h21e0 : data <= 32'h2320f4fe;
	16'h21e1 : data <= 32'h832704fe;
	16'h21e2 : data <= 32'h93f707fc;
	16'h21e3 : data <= 32'h2320f4fe;
	16'h21e4 : data <= 32'h8327c4fc;
	16'h21e5 : data <= 32'h83a70700;
	16'h21e6 : data <= 32'h032744fc;
	16'h21e7 : data <= 32'h13172700;
	16'h21e8 : data <= 32'h9376f70f;
	16'h21e9 : data <= 32'h032704fe;
	16'h21ea : data <= 32'h33e7e600;
	16'h21eb : data <= 32'h23a2e700;
	16'h21ec : data <= 32'h8327c4fc;
	16'h21ed : data <= 32'h83a70700;
	16'h21ee : data <= 32'h83a74700;
	16'h21ef : data <= 32'h232ef4fc;
	16'h21f0 : data <= 32'h8327c4fd;
	16'h21f1 : data <= 32'h93f7e7ff;
	16'h21f2 : data <= 32'h232ef4fc;
	16'h21f3 : data <= 32'h8327c4fc;
	16'h21f4 : data <= 32'h83a70700;
	16'h21f5 : data <= 32'h0327c4fd;
	16'h21f6 : data <= 32'h23a2e700;
	16'h21f7 : data <= 32'h8327c4fc;
	16'h21f8 : data <= 32'h83a70700;
	16'h21f9 : data <= 32'h83a74700;
	16'h21fa : data <= 32'h232cf4fc;
	16'h21fb : data <= 32'h832784fd;
	16'h21fc : data <= 32'h93f7e7ff;
	16'h21fd : data <= 32'h232cf4fc;
	16'h21fe : data <= 32'h8327c4fc;
	16'h21ff : data <= 32'h83a70700;
	16'h2200 : data <= 32'h032784fd;
	16'h2201 : data <= 32'h23a2e700;
	16'h2202 : data <= 32'h6f004001;
	16'h2203 : data <= 32'h8327c4fc;
	16'h2204 : data <= 32'h83a70700;
	16'h2205 : data <= 32'h83a7c700;
	16'h2206 : data <= 32'h232af4fc;
	16'h2207 : data <= 32'h8327c4fc;
	16'h2208 : data <= 32'h83a70700;
	16'h2209 : data <= 32'h83a70701;
	16'h220a : data <= 32'h93d77700;
	16'h220b : data <= 32'h93f71700;
	16'h220c : data <= 32'he38e07fc;
	16'h220d : data <= 32'h8327c4fc;
	16'h220e : data <= 32'h83a70700;
	16'h220f : data <= 32'h83a74700;
	16'h2210 : data <= 32'h2328f4fc;
	16'h2211 : data <= 32'h832704fd;
	16'h2212 : data <= 32'h93f7e7ff;
	16'h2213 : data <= 32'h2328f4fc;
	16'h2214 : data <= 32'h8327c4fc;
	16'h2215 : data <= 32'h83a70700;
	16'h2216 : data <= 32'h032704fd;
	16'h2217 : data <= 32'h13670720;
	16'h2218 : data <= 32'h23a2e700;
	16'h2219 : data <= 32'h8327c4fc;
	16'h221a : data <= 32'h83a70700;
	16'h221b : data <= 32'h83a70701;
	16'h221c : data <= 32'h2324f4fe;
	16'h221d : data <= 32'h6f004008;
	16'h221e : data <= 32'h832784fe;
	16'h221f : data <= 32'h93f71700;
	16'h2220 : data <= 32'h63860700;
	16'h2221 : data <= 32'h93071003;
	16'h2222 : data <= 32'h6f000009;
	16'h2223 : data <= 32'h832784fe;
	16'h2224 : data <= 32'h93d73700;
	16'h2225 : data <= 32'h93f71700;
	16'h2226 : data <= 32'h63860700;
	16'h2227 : data <= 32'h93072003;
	16'h2228 : data <= 32'h6f008007;
	16'h2229 : data <= 32'h832784fe;
	16'h222a : data <= 32'h93d77700;
	16'h222b : data <= 32'h93f71700;
	16'h222c : data <= 32'h639c0702;
	16'h222d : data <= 32'h0327c4fe;
	16'h222e : data <= 32'h832744fc;
	16'h222f : data <= 32'h6376f702;
	16'h2230 : data <= 32'h8327c4fe;
	16'h2231 : data <= 32'h13871700;
	16'h2232 : data <= 32'h2326e4fe;
	16'h2233 : data <= 32'h032784fc;
	16'h2234 : data <= 32'hb307f700;
	16'h2235 : data <= 32'h0327c4fc;
	16'h2236 : data <= 32'h03270700;
	16'h2237 : data <= 32'h0327c700;
	16'h2238 : data <= 32'h1377f70f;
	16'h2239 : data <= 32'h2380e700;
	16'h223a : data <= 32'h8327c4fc;
	16'h223b : data <= 32'h83a70700;
	16'h223c : data <= 32'h83a70701;
	16'h223d : data <= 32'h2324f4fe;
	16'h223e : data <= 32'h0327c4fe;
	16'h223f : data <= 32'h832744fc;
	16'h2240 : data <= 32'he36cf7f6;
	16'h2241 : data <= 32'h832784fe;
	16'h2242 : data <= 32'h93d72700;
	16'h2243 : data <= 32'h93f71700;
	16'h2244 : data <= 32'he38407f6;
	16'h2245 : data <= 32'h93070000;
	16'h2246 : data <= 32'h13850700;
	16'h2247 : data <= 32'h0324c103;
	16'h2248 : data <= 32'h13010104;
	16'h2249 : data <= 32'h67800000;
	16'h224a : data <= 32'h130101fc;
	16'h224b : data <= 32'h232e8102;
	16'h224c : data <= 32'h13040104;
	16'h224d : data <= 32'h2326a4fc;
	16'h224e : data <= 32'h2324b4fc;
	16'h224f : data <= 32'h2322c4fc;
	16'h2250 : data <= 32'h2320d4fc;
	16'h2251 : data <= 32'h232604fe;
	16'h2252 : data <= 32'h032744fc;
	16'h2253 : data <= 32'h93070004;
	16'h2254 : data <= 32'h63f6e700;
	16'h2255 : data <= 32'h93070003;
	16'h2256 : data <= 32'h6f00801d;
	16'h2257 : data <= 32'h032744fc;
	16'h2258 : data <= 32'h93070004;
	16'h2259 : data <= 32'h631af702;
	16'h225a : data <= 32'h8327c4fc;
	16'h225b : data <= 32'h83a70700;
	16'h225c : data <= 32'h83a74700;
	16'h225d : data <= 32'h2324f4fe;
	16'h225e : data <= 32'h832784fe;
	16'h225f : data <= 32'h93f707fc;
	16'h2260 : data <= 32'h2324f4fe;
	16'h2261 : data <= 32'h8327c4fc;
	16'h2262 : data <= 32'h83a70700;
	16'h2263 : data <= 32'h032784fe;
	16'h2264 : data <= 32'h23a2e700;
	16'h2265 : data <= 32'h6f000004;
	16'h2266 : data <= 32'h8327c4fc;
	16'h2267 : data <= 32'h83a70700;
	16'h2268 : data <= 32'h83a74700;
	16'h2269 : data <= 32'h2322f4fe;
	16'h226a : data <= 32'h832744fe;
	16'h226b : data <= 32'h93f707fc;
	16'h226c : data <= 32'h2322f4fe;
	16'h226d : data <= 32'h8327c4fc;
	16'h226e : data <= 32'h83a70700;
	16'h226f : data <= 32'h032744fc;
	16'h2270 : data <= 32'h13172700;
	16'h2271 : data <= 32'h9376f70f;
	16'h2272 : data <= 32'h032744fe;
	16'h2273 : data <= 32'h33e7e600;
	16'h2274 : data <= 32'h23a2e700;
	16'h2275 : data <= 32'h8327c4fc;
	16'h2276 : data <= 32'h83a70700;
	16'h2277 : data <= 32'h83a74700;
	16'h2278 : data <= 32'h2320f4fe;
	16'h2279 : data <= 32'h832704fe;
	16'h227a : data <= 32'h93f7e7ff;
	16'h227b : data <= 32'h2320f4fe;
	16'h227c : data <= 32'h8327c4fc;
	16'h227d : data <= 32'h83a70700;
	16'h227e : data <= 32'h032704fe;
	16'h227f : data <= 32'h13670710;
	16'h2280 : data <= 32'h23a2e700;
	16'h2281 : data <= 32'h8327c4fc;
	16'h2282 : data <= 32'h83a70700;
	16'h2283 : data <= 32'h83a74700;
	16'h2284 : data <= 32'h232ef4fc;
	16'h2285 : data <= 32'h8327c4fd;
	16'h2286 : data <= 32'h93f7e7ff;
	16'h2287 : data <= 32'h232ef4fc;
	16'h2288 : data <= 32'h8327c4fc;
	16'h2289 : data <= 32'h83a70700;
	16'h228a : data <= 32'h0327c4fd;
	16'h228b : data <= 32'h23a2e700;
	16'h228c : data <= 32'h6f000003;
	16'h228d : data <= 32'h8327c4fc;
	16'h228e : data <= 32'h83a70700;
	16'h228f : data <= 32'h032784fc;
	16'h2290 : data <= 32'h03470700;
	16'h2291 : data <= 32'h23a0e700;
	16'h2292 : data <= 32'h832784fc;
	16'h2293 : data <= 32'h93871700;
	16'h2294 : data <= 32'h2324f4fc;
	16'h2295 : data <= 32'h832744fc;
	16'h2296 : data <= 32'h9387f7ff;
	16'h2297 : data <= 32'h2322f4fc;
	16'h2298 : data <= 32'h832744fc;
	16'h2299 : data <= 32'h638e0700;
	16'h229a : data <= 32'h8327c4fc;
	16'h229b : data <= 32'h83a70700;
	16'h229c : data <= 32'h83a70701;
	16'h229d : data <= 32'h93d7b700;
	16'h229e : data <= 32'h93f71700;
	16'h229f : data <= 32'he38c07fa;
	16'h22a0 : data <= 32'h8327c4fc;
	16'h22a1 : data <= 32'h032784fc;
	16'h22a2 : data <= 32'h23a2e700;
	16'h22a3 : data <= 32'h8327c4fc;
	16'h22a4 : data <= 32'h032744fc;
	16'h22a5 : data <= 32'h23a4e700;
	16'h22a6 : data <= 32'h8327c4fc;
	16'h22a7 : data <= 32'h032704fc;
	16'h22a8 : data <= 32'h23a6e700;
	16'h22a9 : data <= 32'h6f008002;
	16'h22aa : data <= 32'h8327c4fc;
	16'h22ab : data <= 32'h03a70700;
	16'h22ac : data <= 32'h8327c4fe;
	16'h22ad : data <= 32'h93861700;
	16'h22ae : data <= 32'h2326d4fe;
	16'h22af : data <= 32'h832684fc;
	16'h22b0 : data <= 32'hb387f600;
	16'h22b1 : data <= 32'h83c70700;
	16'h22b2 : data <= 32'h2320f700;
	16'h22b3 : data <= 32'h0327c4fe;
	16'h22b4 : data <= 32'h832744fc;
	16'h22b5 : data <= 32'h637ef700;
	16'h22b6 : data <= 32'h8327c4fc;
	16'h22b7 : data <= 32'h83a70700;
	16'h22b8 : data <= 32'h83a70701;
	16'h22b9 : data <= 32'h93d7b700;
	16'h22ba : data <= 32'h93f71700;
	16'h22bb : data <= 32'he38e07fa;
	16'h22bc : data <= 32'h8327c4fc;
	16'h22bd : data <= 32'h83a70700;
	16'h22be : data <= 32'h83a74700;
	16'h22bf : data <= 32'h232cf4fc;
	16'h22c0 : data <= 32'h832784fd;
	16'h22c1 : data <= 32'h93f7e7ff;
	16'h22c2 : data <= 32'h232cf4fc;
	16'h22c3 : data <= 32'h8327c4fc;
	16'h22c4 : data <= 32'h83a70700;
	16'h22c5 : data <= 32'h032784fd;
	16'h22c6 : data <= 32'h13670720;
	16'h22c7 : data <= 32'h23a2e700;
	16'h22c8 : data <= 32'h8327c4fc;
	16'h22c9 : data <= 32'h13071000;
	16'h22ca : data <= 32'h23a8e700;
	16'h22cb : data <= 32'h93070000;
	16'h22cc : data <= 32'h13850700;
	16'h22cd : data <= 32'h0324c103;
	16'h22ce : data <= 32'h13010104;
	16'h22cf : data <= 32'h67800000;
	16'h22d0 : data <= 32'h130101fd;
	16'h22d1 : data <= 32'h23268102;
	16'h22d2 : data <= 32'h13040103;
	16'h22d3 : data <= 32'h232ea4fc;
	16'h22d4 : data <= 32'h232cb4fc;
	16'h22d5 : data <= 32'h232ac4fc;
	16'h22d6 : data <= 32'h232604fe;
	16'h22d7 : data <= 32'h8327c4fd;
	16'h22d8 : data <= 32'h83a70700;
	16'h22d9 : data <= 32'h83a74700;
	16'h22da : data <= 32'h2322f4fe;
	16'h22db : data <= 32'h832744fe;
	16'h22dc : data <= 32'h93f7e7ff;
	16'h22dd : data <= 32'h2322f4fe;
	16'h22de : data <= 32'h8327c4fd;
	16'h22df : data <= 32'h83a70700;
	16'h22e0 : data <= 32'h032744fe;
	16'h22e1 : data <= 32'h13672700;
	16'h22e2 : data <= 32'h23a2e700;
	16'h22e3 : data <= 32'h6f008002;
	16'h22e4 : data <= 32'h8327c4fd;
	16'h22e5 : data <= 32'h03a70700;
	16'h22e6 : data <= 32'h8327c4fe;
	16'h22e7 : data <= 32'h93861700;
	16'h22e8 : data <= 32'h2326d4fe;
	16'h22e9 : data <= 32'h832684fd;
	16'h22ea : data <= 32'hb387f600;
	16'h22eb : data <= 32'h83c70700;
	16'h22ec : data <= 32'h2320f700;
	16'h22ed : data <= 32'h0327c4fe;
	16'h22ee : data <= 32'h832744fd;
	16'h22ef : data <= 32'h637ef700;
	16'h22f0 : data <= 32'h8327c4fd;
	16'h22f1 : data <= 32'h83a70700;
	16'h22f2 : data <= 32'h83a70701;
	16'h22f3 : data <= 32'h93d7b700;
	16'h22f4 : data <= 32'h93f71700;
	16'h22f5 : data <= 32'he38e07fa;
	16'h22f6 : data <= 32'h8327c4fd;
	16'h22f7 : data <= 32'h83a70700;
	16'h22f8 : data <= 32'h83a70701;
	16'h22f9 : data <= 32'h2324f4fe;
	16'h22fa : data <= 32'h6f008006;
	16'h22fb : data <= 32'h832784fe;
	16'h22fc : data <= 32'h93f71700;
	16'h22fd : data <= 32'h63860700;
	16'h22fe : data <= 32'h93071003;
	16'h22ff : data <= 32'h6f004007;
	16'h2300 : data <= 32'h832784fe;
	16'h2301 : data <= 32'h93d7b700;
	16'h2302 : data <= 32'h93f71700;
	16'h2303 : data <= 32'h639a0702;
	16'h2304 : data <= 32'h0327c4fe;
	16'h2305 : data <= 32'h832744fd;
	16'h2306 : data <= 32'h6374f702;
	16'h2307 : data <= 32'h8327c4fd;
	16'h2308 : data <= 32'h03a70700;
	16'h2309 : data <= 32'h8327c4fe;
	16'h230a : data <= 32'h93861700;
	16'h230b : data <= 32'h2326d4fe;
	16'h230c : data <= 32'h832684fd;
	16'h230d : data <= 32'hb387f600;
	16'h230e : data <= 32'h83c70700;
	16'h230f : data <= 32'h2320f700;
	16'h2310 : data <= 32'h8327c4fd;
	16'h2311 : data <= 32'h83a70700;
	16'h2312 : data <= 32'h83a70701;
	16'h2313 : data <= 32'h2324f4fe;
	16'h2314 : data <= 32'h0327c4fe;
	16'h2315 : data <= 32'h832744fd;
	16'h2316 : data <= 32'he36af7f8;
	16'h2317 : data <= 32'h832784fe;
	16'h2318 : data <= 32'h93d72700;
	16'h2319 : data <= 32'h93f71700;
	16'h231a : data <= 32'he38207f8;
	16'h231b : data <= 32'h93070000;
	16'h231c : data <= 32'h13850700;
	16'h231d : data <= 32'h0324c102;
	16'h231e : data <= 32'h13010103;
	16'h231f : data <= 32'h67800000;
	16'h2320 : data <= 32'h130101fd;
	16'h2321 : data <= 32'h23268102;
	16'h2322 : data <= 32'h13040103;
	16'h2323 : data <= 32'h232ea4fc;
	16'h2324 : data <= 32'h232cb4fc;
	16'h2325 : data <= 32'h232ac4fc;
	16'h2326 : data <= 32'h232604fe;
	16'h2327 : data <= 32'h8327c4fd;
	16'h2328 : data <= 32'h83a70700;
	16'h2329 : data <= 32'h83a74700;
	16'h232a : data <= 32'h2322f4fe;
	16'h232b : data <= 32'h832744fe;
	16'h232c : data <= 32'h93f7e7ff;
	16'h232d : data <= 32'h2322f4fe;
	16'h232e : data <= 32'h8327c4fd;
	16'h232f : data <= 32'h83a70700;
	16'h2330 : data <= 32'h032744fe;
	16'h2331 : data <= 32'h13672700;
	16'h2332 : data <= 32'h23a2e700;
	16'h2333 : data <= 32'h6f004001;
	16'h2334 : data <= 32'h8327c4fd;
	16'h2335 : data <= 32'h83a70700;
	16'h2336 : data <= 32'h83a7c700;
	16'h2337 : data <= 32'h2320f4fe;
	16'h2338 : data <= 32'h8327c4fd;
	16'h2339 : data <= 32'h83a70700;
	16'h233a : data <= 32'h83a70701;
	16'h233b : data <= 32'h93d77700;
	16'h233c : data <= 32'h93f71700;
	16'h233d : data <= 32'he38e07fc;
	16'h233e : data <= 32'h8327c4fd;
	16'h233f : data <= 32'h83a70700;
	16'h2340 : data <= 32'h83a70701;
	16'h2341 : data <= 32'h2324f4fe;
	16'h2342 : data <= 32'h6f00c006;
	16'h2343 : data <= 32'h832784fe;
	16'h2344 : data <= 32'h93f71700;
	16'h2345 : data <= 32'h63860700;
	16'h2346 : data <= 32'h93071003;
	16'h2347 : data <= 32'h6f008007;
	16'h2348 : data <= 32'h832784fe;
	16'h2349 : data <= 32'h93d77700;
	16'h234a : data <= 32'h93f71700;
	16'h234b : data <= 32'h639c0702;
	16'h234c : data <= 32'h0327c4fe;
	16'h234d : data <= 32'h832744fd;
	16'h234e : data <= 32'h6376f702;
	16'h234f : data <= 32'h8327c4fe;
	16'h2350 : data <= 32'h13871700;
	16'h2351 : data <= 32'h2326e4fe;
	16'h2352 : data <= 32'h032784fd;
	16'h2353 : data <= 32'hb307f700;
	16'h2354 : data <= 32'h0327c4fd;
	16'h2355 : data <= 32'h03270700;
	16'h2356 : data <= 32'h0327c700;
	16'h2357 : data <= 32'h1377f70f;
	16'h2358 : data <= 32'h2380e700;
	16'h2359 : data <= 32'h8327c4fd;
	16'h235a : data <= 32'h83a70700;
	16'h235b : data <= 32'h83a70701;
	16'h235c : data <= 32'h2324f4fe;
	16'h235d : data <= 32'h0327c4fe;
	16'h235e : data <= 32'h832744fd;
	16'h235f : data <= 32'he368f7f8;
	16'h2360 : data <= 32'h832784fe;
	16'h2361 : data <= 32'h93d72700;
	16'h2362 : data <= 32'h93f71700;
	16'h2363 : data <= 32'he38007f8;
	16'h2364 : data <= 32'h93070000;
	16'h2365 : data <= 32'h13850700;
	16'h2366 : data <= 32'h0324c102;
	16'h2367 : data <= 32'h13010103;
	16'h2368 : data <= 32'h67800000;
	16'h2369 : data <= 32'h130101fd;
	16'h236a : data <= 32'h23268102;
	16'h236b : data <= 32'h13040103;
	16'h236c : data <= 32'h232ea4fc;
	16'h236d : data <= 32'h232cb4fc;
	16'h236e : data <= 32'h232ac4fc;
	16'h236f : data <= 32'h2328d4fc;
	16'h2370 : data <= 32'h232604fe;
	16'h2371 : data <= 32'h8327c4fd;
	16'h2372 : data <= 32'h83a70700;
	16'h2373 : data <= 32'h83a74700;
	16'h2374 : data <= 32'h2324f4fe;
	16'h2375 : data <= 32'h832784fe;
	16'h2376 : data <= 32'h93f7e7ff;
	16'h2377 : data <= 32'h2324f4fe;
	16'h2378 : data <= 32'h8327c4fd;
	16'h2379 : data <= 32'h83a70700;
	16'h237a : data <= 32'h032784fe;
	16'h237b : data <= 32'h13672700;
	16'h237c : data <= 32'h23a2e700;
	16'h237d : data <= 32'h6f000003;
	16'h237e : data <= 32'h8327c4fd;
	16'h237f : data <= 32'h83a70700;
	16'h2380 : data <= 32'h032784fd;
	16'h2381 : data <= 32'h03470700;
	16'h2382 : data <= 32'h23a0e700;
	16'h2383 : data <= 32'h832784fd;
	16'h2384 : data <= 32'h93871700;
	16'h2385 : data <= 32'h232cf4fc;
	16'h2386 : data <= 32'h832744fd;
	16'h2387 : data <= 32'h9387f7ff;
	16'h2388 : data <= 32'h232af4fc;
	16'h2389 : data <= 32'h832744fd;
	16'h238a : data <= 32'h638e0700;
	16'h238b : data <= 32'h8327c4fd;
	16'h238c : data <= 32'h83a70700;
	16'h238d : data <= 32'h83a70701;
	16'h238e : data <= 32'h93d7b700;
	16'h238f : data <= 32'h93f71700;
	16'h2390 : data <= 32'he38c07fa;
	16'h2391 : data <= 32'h8327c4fd;
	16'h2392 : data <= 32'h032784fd;
	16'h2393 : data <= 32'h23a2e700;
	16'h2394 : data <= 32'h8327c4fd;
	16'h2395 : data <= 32'h032744fd;
	16'h2396 : data <= 32'h23a4e700;
	16'h2397 : data <= 32'h8327c4fd;
	16'h2398 : data <= 32'h032704fd;
	16'h2399 : data <= 32'h23a6e700;
	16'h239a : data <= 32'h6f008002;
	16'h239b : data <= 32'h8327c4fd;
	16'h239c : data <= 32'h03a70700;
	16'h239d : data <= 32'h8327c4fe;
	16'h239e : data <= 32'h93861700;
	16'h239f : data <= 32'h2326d4fe;
	16'h23a0 : data <= 32'h832684fd;
	16'h23a1 : data <= 32'hb387f600;
	16'h23a2 : data <= 32'h83c70700;
	16'h23a3 : data <= 32'h2320f700;
	16'h23a4 : data <= 32'h0327c4fe;
	16'h23a5 : data <= 32'h832744fd;
	16'h23a6 : data <= 32'h637ef700;
	16'h23a7 : data <= 32'h8327c4fd;
	16'h23a8 : data <= 32'h83a70700;
	16'h23a9 : data <= 32'h83a70701;
	16'h23aa : data <= 32'h93d7b700;
	16'h23ab : data <= 32'h93f71700;
	16'h23ac : data <= 32'he38e07fa;
	16'h23ad : data <= 32'h8327c4fd;
	16'h23ae : data <= 32'h13071000;
	16'h23af : data <= 32'h23a8e700;
	16'h23b0 : data <= 32'h93070000;
	16'h23b1 : data <= 32'h13850700;
	16'h23b2 : data <= 32'h0324c102;
	16'h23b3 : data <= 32'h13010103;
	16'h23b4 : data <= 32'h67800000;
	16'h23b5 : data <= 32'h130101fd;
	16'h23b6 : data <= 32'h23268102;
	16'h23b7 : data <= 32'h13040103;
	16'h23b8 : data <= 32'h232ea4fc;
	16'h23b9 : data <= 32'h232cb4fc;
	16'h23ba : data <= 32'h232ac4fc;
	16'h23bb : data <= 32'h2328d4fc;
	16'h23bc : data <= 32'h232604fe;
	16'h23bd : data <= 32'h8327c4fd;
	16'h23be : data <= 32'h83a70700;
	16'h23bf : data <= 32'h83a74700;
	16'h23c0 : data <= 32'h2324f4fe;
	16'h23c1 : data <= 32'h832784fe;
	16'h23c2 : data <= 32'h93f7e7ff;
	16'h23c3 : data <= 32'h2324f4fe;
	16'h23c4 : data <= 32'h8327c4fd;
	16'h23c5 : data <= 32'h83a70700;
	16'h23c6 : data <= 32'h032784fe;
	16'h23c7 : data <= 32'h13672700;
	16'h23c8 : data <= 32'h23a2e700;
	16'h23c9 : data <= 32'h6f004001;
	16'h23ca : data <= 32'h8327c4fd;
	16'h23cb : data <= 32'h83a70700;
	16'h23cc : data <= 32'h83a7c700;
	16'h23cd : data <= 32'h2322f4fe;
	16'h23ce : data <= 32'h8327c4fd;
	16'h23cf : data <= 32'h83a70700;
	16'h23d0 : data <= 32'h83a70701;
	16'h23d1 : data <= 32'h93d77700;
	16'h23d2 : data <= 32'h93f71700;
	16'h23d3 : data <= 32'he38e07fc;
	16'h23d4 : data <= 32'h8327c4fd;
	16'h23d5 : data <= 32'h032784fd;
	16'h23d6 : data <= 32'h23a2e700;
	16'h23d7 : data <= 32'h8327c4fd;
	16'h23d8 : data <= 32'h032744fd;
	16'h23d9 : data <= 32'h23a4e700;
	16'h23da : data <= 32'h8327c4fd;
	16'h23db : data <= 32'h032704fd;
	16'h23dc : data <= 32'h23a6e700;
	16'h23dd : data <= 32'h8327c4fd;
	16'h23de : data <= 32'h13072000;
	16'h23df : data <= 32'h23a8e700;
	16'h23e0 : data <= 32'h93070000;
	16'h23e1 : data <= 32'h13850700;
	16'h23e2 : data <= 32'h0324c102;
	16'h23e3 : data <= 32'h13010103;
	16'h23e4 : data <= 32'h67800000;
	16'h23e5 : data <= 32'h130101fd;
	16'h23e6 : data <= 32'h23261102;
	16'h23e7 : data <= 32'h23248102;
	16'h23e8 : data <= 32'h13040103;
	16'h23e9 : data <= 32'h232ea4fc;
	16'h23ea : data <= 32'h8327c4fd;
	16'h23eb : data <= 32'h03a70701;
	16'h23ec : data <= 32'h93071000;
	16'h23ed : data <= 32'h630af700;
	16'h23ee : data <= 32'h8327c4fd;
	16'h23ef : data <= 32'h03a70701;
	16'h23f0 : data <= 32'h93072000;
	16'h23f1 : data <= 32'h631cf718;
	16'h23f2 : data <= 32'h8327c4fd;
	16'h23f3 : data <= 32'h83a70700;
	16'h23f4 : data <= 32'h83a70701;
	16'h23f5 : data <= 32'h2326f4fe;
	16'h23f6 : data <= 32'h8327c4fe;
	16'h23f7 : data <= 32'h93f71700;
	16'h23f8 : data <= 32'h63820702;
	16'h23f9 : data <= 32'h8327c4fd;
	16'h23fa : data <= 32'h13073000;
	16'h23fb : data <= 32'h23a8e700;
	16'h23fc : data <= 32'h8327c4fd;
	16'h23fd : data <= 32'h83a7c700;
	16'h23fe : data <= 32'h13051003;
	16'h23ff : data <= 32'he7800700;
	16'h2400 : data <= 32'h6f000016;
	16'h2401 : data <= 32'h8327c4fe;
	16'h2402 : data <= 32'h93d73700;
	16'h2403 : data <= 32'h93f71700;
	16'h2404 : data <= 32'h63820702;
	16'h2405 : data <= 32'h8327c4fd;
	16'h2406 : data <= 32'h13073000;
	16'h2407 : data <= 32'h23a8e700;
	16'h2408 : data <= 32'h8327c4fd;
	16'h2409 : data <= 32'h83a7c700;
	16'h240a : data <= 32'h13052003;
	16'h240b : data <= 32'he7800700;
	16'h240c : data <= 32'h6f000013;
	16'h240d : data <= 32'h8327c4fe;
	16'h240e : data <= 32'h93d72700;
	16'h240f : data <= 32'h93f71700;
	16'h2410 : data <= 32'h63820702;
	16'h2411 : data <= 32'h8327c4fd;
	16'h2412 : data <= 32'h13073000;
	16'h2413 : data <= 32'h23a8e700;
	16'h2414 : data <= 32'h8327c4fd;
	16'h2415 : data <= 32'h83a7c700;
	16'h2416 : data <= 32'h13050000;
	16'h2417 : data <= 32'he7800700;
	16'h2418 : data <= 32'h6f000010;
	16'h2419 : data <= 32'h8327c4fd;
	16'h241a : data <= 32'h03a70701;
	16'h241b : data <= 32'h93071000;
	16'h241c : data <= 32'h6316f70c;
	16'h241d : data <= 32'h6f004005;
	16'h241e : data <= 32'h8327c4fd;
	16'h241f : data <= 32'h83a70700;
	16'h2420 : data <= 32'h0327c4fd;
	16'h2421 : data <= 32'h03274700;
	16'h2422 : data <= 32'h03470700;
	16'h2423 : data <= 32'h23a0e700;
	16'h2424 : data <= 32'h8327c4fd;
	16'h2425 : data <= 32'h83a74700;
	16'h2426 : data <= 32'h13871700;
	16'h2427 : data <= 32'h8327c4fd;
	16'h2428 : data <= 32'h23a2e700;
	16'h2429 : data <= 32'h8327c4fd;
	16'h242a : data <= 32'h83a78700;
	16'h242b : data <= 32'h1387f7ff;
	16'h242c : data <= 32'h8327c4fd;
	16'h242d : data <= 32'h23a4e700;
	16'h242e : data <= 32'h8327c4fd;
	16'h242f : data <= 32'h83a70700;
	16'h2430 : data <= 32'h83a70701;
	16'h2431 : data <= 32'h2326f4fe;
	16'h2432 : data <= 32'h8327c4fe;
	16'h2433 : data <= 32'h93d7b700;
	16'h2434 : data <= 32'h93f71700;
	16'h2435 : data <= 32'h63960708;
	16'h2436 : data <= 32'h8327c4fd;
	16'h2437 : data <= 32'h83a78700;
	16'h2438 : data <= 32'he39c07f8;
	16'h2439 : data <= 32'h6f00c007;
	16'h243a : data <= 32'h8327c4fd;
	16'h243b : data <= 32'h83a74700;
	16'h243c : data <= 32'h0327c4fd;
	16'h243d : data <= 32'h03270700;
	16'h243e : data <= 32'h0327c700;
	16'h243f : data <= 32'h1377f70f;
	16'h2440 : data <= 32'h2380e700;
	16'h2441 : data <= 32'h8327c4fd;
	16'h2442 : data <= 32'h83a74700;
	16'h2443 : data <= 32'h13871700;
	16'h2444 : data <= 32'h8327c4fd;
	16'h2445 : data <= 32'h23a2e700;
	16'h2446 : data <= 32'h8327c4fd;
	16'h2447 : data <= 32'h83a78700;
	16'h2448 : data <= 32'h1387f7ff;
	16'h2449 : data <= 32'h8327c4fd;
	16'h244a : data <= 32'h23a4e700;
	16'h244b : data <= 32'h8327c4fd;
	16'h244c : data <= 32'h83a70700;
	16'h244d : data <= 32'h83a70701;
	16'h244e : data <= 32'h2326f4fe;
	16'h244f : data <= 32'h8327c4fe;
	16'h2450 : data <= 32'h93d77700;
	16'h2451 : data <= 32'h93f71700;
	16'h2452 : data <= 32'h639c0700;
	16'h2453 : data <= 32'h8327c4fd;
	16'h2454 : data <= 32'h83a78700;
	16'h2455 : data <= 32'he39a07f8;
	16'h2456 : data <= 32'h6f008000;
	16'h2457 : data <= 32'h13000000;
	16'h2458 : data <= 32'h8320c102;
	16'h2459 : data <= 32'h03248102;
	16'h245a : data <= 32'h13010103;
	16'h245b : data <= 32'h67800000;
	16'h245c : data <= 32'h130101fc;
	16'h245d : data <= 32'h232e8102;
	16'h245e : data <= 32'h13040104;
	16'h245f : data <= 32'h2326a4fc;
	16'h2460 : data <= 32'h2324b4fc;
	16'h2461 : data <= 32'h2322c4fc;
	16'h2462 : data <= 32'h2320d4fc;
	16'h2463 : data <= 32'h232604fe;
	16'h2464 : data <= 32'h032744fc;
	16'h2465 : data <= 32'h93070004;
	16'h2466 : data <= 32'h63f6e700;
	16'h2467 : data <= 32'h93070003;
	16'h2468 : data <= 32'h6f004016;
	16'h2469 : data <= 32'h032744fc;
	16'h246a : data <= 32'h93070004;
	16'h246b : data <= 32'h631af702;
	16'h246c : data <= 32'h8327c4fc;
	16'h246d : data <= 32'h83a70700;
	16'h246e : data <= 32'h83a74700;
	16'h246f : data <= 32'h2324f4fe;
	16'h2470 : data <= 32'h832784fe;
	16'h2471 : data <= 32'h93f707fc;
	16'h2472 : data <= 32'h2324f4fe;
	16'h2473 : data <= 32'h8327c4fc;
	16'h2474 : data <= 32'h83a70700;
	16'h2475 : data <= 32'h032784fe;
	16'h2476 : data <= 32'h23a2e700;
	16'h2477 : data <= 32'h6f000004;
	16'h2478 : data <= 32'h8327c4fc;
	16'h2479 : data <= 32'h83a70700;
	16'h247a : data <= 32'h83a74700;
	16'h247b : data <= 32'h2322f4fe;
	16'h247c : data <= 32'h832744fe;
	16'h247d : data <= 32'h93f707fc;
	16'h247e : data <= 32'h2322f4fe;
	16'h247f : data <= 32'h8327c4fc;
	16'h2480 : data <= 32'h83a70700;
	16'h2481 : data <= 32'h032744fc;
	16'h2482 : data <= 32'h13172700;
	16'h2483 : data <= 32'h9376f70f;
	16'h2484 : data <= 32'h032744fe;
	16'h2485 : data <= 32'h33e7e600;
	16'h2486 : data <= 32'h23a2e700;
	16'h2487 : data <= 32'h8327c4fc;
	16'h2488 : data <= 32'h83a70700;
	16'h2489 : data <= 32'h83a74700;
	16'h248a : data <= 32'h2320f4fe;
	16'h248b : data <= 32'h832704fe;
	16'h248c : data <= 32'h93f7e7ff;
	16'h248d : data <= 32'h2320f4fe;
	16'h248e : data <= 32'h8327c4fc;
	16'h248f : data <= 32'h83a70700;
	16'h2490 : data <= 32'h032704fe;
	16'h2491 : data <= 32'h23a2e700;
	16'h2492 : data <= 32'h8327c4fc;
	16'h2493 : data <= 32'h83a70700;
	16'h2494 : data <= 32'h83a74700;
	16'h2495 : data <= 32'h232ef4fc;
	16'h2496 : data <= 32'h8327c4fd;
	16'h2497 : data <= 32'h93f7e7ff;
	16'h2498 : data <= 32'h232ef4fc;
	16'h2499 : data <= 32'h8327c4fc;
	16'h249a : data <= 32'h83a70700;
	16'h249b : data <= 32'h0327c4fd;
	16'h249c : data <= 32'h23a2e700;
	16'h249d : data <= 32'h6f004001;
	16'h249e : data <= 32'h8327c4fc;
	16'h249f : data <= 32'h83a70700;
	16'h24a0 : data <= 32'h83a7c700;
	16'h24a1 : data <= 32'h232cf4fc;
	16'h24a2 : data <= 32'h8327c4fc;
	16'h24a3 : data <= 32'h83a70700;
	16'h24a4 : data <= 32'h83a70701;
	16'h24a5 : data <= 32'h93d77700;
	16'h24a6 : data <= 32'h93f71700;
	16'h24a7 : data <= 32'he38e07fc;
	16'h24a8 : data <= 32'h8327c4fc;
	16'h24a9 : data <= 32'h032784fc;
	16'h24aa : data <= 32'h23a2e700;
	16'h24ab : data <= 32'h8327c4fc;
	16'h24ac : data <= 32'h032744fc;
	16'h24ad : data <= 32'h23a4e700;
	16'h24ae : data <= 32'h8327c4fc;
	16'h24af : data <= 32'h032704fc;
	16'h24b0 : data <= 32'h23a6e700;
	16'h24b1 : data <= 32'h8327c4fc;
	16'h24b2 : data <= 32'h83a70700;
	16'h24b3 : data <= 32'h83a74700;
	16'h24b4 : data <= 32'h232af4fc;
	16'h24b5 : data <= 32'h832744fd;
	16'h24b6 : data <= 32'h93f7e7ff;
	16'h24b7 : data <= 32'h232af4fc;
	16'h24b8 : data <= 32'h8327c4fc;
	16'h24b9 : data <= 32'h83a70700;
	16'h24ba : data <= 32'h032744fd;
	16'h24bb : data <= 32'h13670720;
	16'h24bc : data <= 32'h23a2e700;
	16'h24bd : data <= 32'h8327c4fc;
	16'h24be : data <= 32'h13072000;
	16'h24bf : data <= 32'h23a8e700;
	16'h24c0 : data <= 32'h93070000;
	16'h24c1 : data <= 32'h13850700;
	16'h24c2 : data <= 32'h0324c103;
	16'h24c3 : data <= 32'h13010104;
	16'h24c4 : data <= 32'h67800000;
	16'h24c5 : data <= 32'h130101fd;
	16'h24c6 : data <= 32'h23268102;
	16'h24c7 : data <= 32'h13040103;
	16'h24c8 : data <= 32'h232ea4fc;
	16'h24c9 : data <= 32'h232cb4fc;
	16'h24ca : data <= 32'h232ac4fc;
	16'h24cb : data <= 32'h232604fe;
	16'h24cc : data <= 32'h232604fe;
	16'h24cd : data <= 32'h6f008004;
	16'h24ce : data <= 32'h13000000;
	16'h24cf : data <= 32'h8327c4fd;
	16'h24d0 : data <= 32'h83a70700;
	16'h24d1 : data <= 32'h83a7c700;
	16'h24d2 : data <= 32'h93d72700;
	16'h24d3 : data <= 32'h93f71700;
	16'h24d4 : data <= 32'he39607fe;
	16'h24d5 : data <= 32'h8327c4fd;
	16'h24d6 : data <= 32'h83a70700;
	16'h24d7 : data <= 32'h0327c4fe;
	16'h24d8 : data <= 32'h832684fd;
	16'h24d9 : data <= 32'h3387e600;
	16'h24da : data <= 32'h03470700;
	16'h24db : data <= 32'h23a2e700;
	16'h24dc : data <= 32'h8327c4fe;
	16'h24dd : data <= 32'h93871700;
	16'h24de : data <= 32'h2326f4fe;
	16'h24df : data <= 32'h0327c4fe;
	16'h24e0 : data <= 32'h832744fd;
	16'h24e1 : data <= 32'he36af7fa;
	16'h24e2 : data <= 32'h93070000;
	16'h24e3 : data <= 32'h13850700;
	16'h24e4 : data <= 32'h0324c102;
	16'h24e5 : data <= 32'h13010103;
	16'h24e6 : data <= 32'h67800000;
	16'h24e7 : data <= 32'h130101fd;
	16'h24e8 : data <= 32'h23268102;
	16'h24e9 : data <= 32'h13040103;
	16'h24ea : data <= 32'h232ea4fc;
	16'h24eb : data <= 32'h232cb4fc;
	16'h24ec : data <= 32'h232ac4fc;
	16'h24ed : data <= 32'h232604fe;
	16'h24ee : data <= 32'h232604fe;
	16'h24ef : data <= 32'h6f00c004;
	16'h24f0 : data <= 32'h13000000;
	16'h24f1 : data <= 32'h8327c4fd;
	16'h24f2 : data <= 32'h83a70700;
	16'h24f3 : data <= 32'h83a7c700;
	16'h24f4 : data <= 32'h93d75700;
	16'h24f5 : data <= 32'h93f71700;
	16'h24f6 : data <= 32'he39607fe;
	16'h24f7 : data <= 32'h8327c4fe;
	16'h24f8 : data <= 32'h032784fd;
	16'h24f9 : data <= 32'hb307f700;
	16'h24fa : data <= 32'h0327c4fd;
	16'h24fb : data <= 32'h03270700;
	16'h24fc : data <= 32'h03278700;
	16'h24fd : data <= 32'h1377f70f;
	16'h24fe : data <= 32'h2380e700;
	16'h24ff : data <= 32'h8327c4fe;
	16'h2500 : data <= 32'h93871700;
	16'h2501 : data <= 32'h2326f4fe;
	16'h2502 : data <= 32'h0327c4fe;
	16'h2503 : data <= 32'h832744fd;
	16'h2504 : data <= 32'he368f7fa;
	16'h2505 : data <= 32'h93070000;
	16'h2506 : data <= 32'h13850700;
	16'h2507 : data <= 32'h0324c102;
	16'h2508 : data <= 32'h13010103;
	16'h2509 : data <= 32'h67800000;
	16'h250a : data <= 32'h130101fe;
	16'h250b : data <= 32'h232e1100;
	16'h250c : data <= 32'h232c8100;
	16'h250d : data <= 32'h13040102;
	16'h250e : data <= 32'h2326a4fe;
	16'h250f : data <= 32'h2324b4fe;
	16'h2510 : data <= 32'h2322c4fe;
	16'h2511 : data <= 32'h2320d4fe;
	16'h2512 : data <= 32'h8327c4fe;
	16'h2513 : data <= 32'h83a70702;
	16'h2514 : data <= 32'h63960700;
	16'h2515 : data <= 32'h93070002;
	16'h2516 : data <= 32'h6f00c00c;
	16'h2517 : data <= 32'h8327c4fe;
	16'h2518 : data <= 32'h03a70702;
	16'h2519 : data <= 32'h93071000;
	16'h251a : data <= 32'h6316f700;
	16'h251b : data <= 32'h93071002;
	16'h251c : data <= 32'h6f00400b;
	16'h251d : data <= 32'h8327c4fe;
	16'h251e : data <= 32'h03a70702;
	16'h251f : data <= 32'h93072000;
	16'h2520 : data <= 32'h630cf702;
	16'h2521 : data <= 32'h93071000;
	16'h2522 : data <= 32'h6f00c009;
	16'h2523 : data <= 32'h8327c4fe;
	16'h2524 : data <= 32'h83a70700;
	16'h2525 : data <= 32'h032784fe;
	16'h2526 : data <= 32'h03470700;
	16'h2527 : data <= 32'h23a2e700;
	16'h2528 : data <= 32'h832784fe;
	16'h2529 : data <= 32'h93871700;
	16'h252a : data <= 32'h2324f4fe;
	16'h252b : data <= 32'h832744fe;
	16'h252c : data <= 32'h9387f7ff;
	16'h252d : data <= 32'h2322f4fe;
	16'h252e : data <= 32'h832744fe;
	16'h252f : data <= 32'h638e0700;
	16'h2530 : data <= 32'h8327c4fe;
	16'h2531 : data <= 32'h83a70700;
	16'h2532 : data <= 32'h83a7c700;
	16'h2533 : data <= 32'h93d72700;
	16'h2534 : data <= 32'h93f71700;
	16'h2535 : data <= 32'he38c07fa;
	16'h2536 : data <= 32'h832744fe;
	16'h2537 : data <= 32'h639a0700;
	16'h2538 : data <= 32'h832704fe;
	16'h2539 : data <= 32'he7800700;
	16'h253a : data <= 32'h93070000;
	16'h253b : data <= 32'h6f008003;
	16'h253c : data <= 32'h8327c4fe;
	16'h253d : data <= 32'h032784fe;
	16'h253e : data <= 32'h23a2e700;
	16'h253f : data <= 32'h8327c4fe;
	16'h2540 : data <= 32'h032744fe;
	16'h2541 : data <= 32'h23a6e700;
	16'h2542 : data <= 32'h8327c4fe;
	16'h2543 : data <= 32'h032704fe;
	16'h2544 : data <= 32'h23aae700;
	16'h2545 : data <= 32'h8327c4fe;
	16'h2546 : data <= 32'h13071000;
	16'h2547 : data <= 32'h23a0e702;
	16'h2548 : data <= 32'h93070000;
	16'h2549 : data <= 32'h13850700;
	16'h254a : data <= 32'h8320c101;
	16'h254b : data <= 32'h03248101;
	16'h254c : data <= 32'h13010102;
	16'h254d : data <= 32'h67800000;
	16'h254e : data <= 32'h130101fe;
	16'h254f : data <= 32'h232e1100;
	16'h2550 : data <= 32'h232c8100;
	16'h2551 : data <= 32'h13040102;
	16'h2552 : data <= 32'h2326a4fe;
	16'h2553 : data <= 32'h2324b4fe;
	16'h2554 : data <= 32'h93070600;
	16'h2555 : data <= 32'h2320d4fe;
	16'h2556 : data <= 32'h2313f4fe;
	16'h2557 : data <= 32'h8327c4fe;
	16'h2558 : data <= 32'h83a70702;
	16'h2559 : data <= 32'h63960700;
	16'h255a : data <= 32'h93070002;
	16'h255b : data <= 32'h6f00000d;
	16'h255c : data <= 32'h8327c4fe;
	16'h255d : data <= 32'h03a70702;
	16'h255e : data <= 32'h93071000;
	16'h255f : data <= 32'h6316f700;
	16'h2560 : data <= 32'h93071002;
	16'h2561 : data <= 32'h6f00800b;
	16'h2562 : data <= 32'h8327c4fe;
	16'h2563 : data <= 32'h03a70702;
	16'h2564 : data <= 32'h93072000;
	16'h2565 : data <= 32'h630ef702;
	16'h2566 : data <= 32'h93071000;
	16'h2567 : data <= 32'h6f00000a;
	16'h2568 : data <= 32'h8327c4fe;
	16'h2569 : data <= 32'h83a70700;
	16'h256a : data <= 32'h83a78700;
	16'h256b : data <= 32'h13f7f70f;
	16'h256c : data <= 32'h832784fe;
	16'h256d : data <= 32'h2380e700;
	16'h256e : data <= 32'h832784fe;
	16'h256f : data <= 32'h93871700;
	16'h2570 : data <= 32'h2324f4fe;
	16'h2571 : data <= 32'h835764fe;
	16'h2572 : data <= 32'h9387f7ff;
	16'h2573 : data <= 32'h2313f4fe;
	16'h2574 : data <= 32'h835764fe;
	16'h2575 : data <= 32'h638e0700;
	16'h2576 : data <= 32'h8327c4fe;
	16'h2577 : data <= 32'h83a70700;
	16'h2578 : data <= 32'h83a7c700;
	16'h2579 : data <= 32'h93d75700;
	16'h257a : data <= 32'h93f71700;
	16'h257b : data <= 32'he38a07fa;
	16'h257c : data <= 32'h835764fe;
	16'h257d : data <= 32'h639a0700;
	16'h257e : data <= 32'h832704fe;
	16'h257f : data <= 32'he7800700;
	16'h2580 : data <= 32'h93070000;
	16'h2581 : data <= 32'h6f008003;
	16'h2582 : data <= 32'h8327c4fe;
	16'h2583 : data <= 32'h032784fe;
	16'h2584 : data <= 32'h23a4e700;
	16'h2585 : data <= 32'h035764fe;
	16'h2586 : data <= 32'h8327c4fe;
	16'h2587 : data <= 32'h23a8e700;
	16'h2588 : data <= 32'h8327c4fe;
	16'h2589 : data <= 32'h032704fe;
	16'h258a : data <= 32'h23ace700;
	16'h258b : data <= 32'h8327c4fe;
	16'h258c : data <= 32'h13071000;
	16'h258d : data <= 32'h23aee700;
	16'h258e : data <= 32'h93070000;
	16'h258f : data <= 32'h13850700;
	16'h2590 : data <= 32'h8320c101;
	16'h2591 : data <= 32'h03248101;
	16'h2592 : data <= 32'h13010102;
	16'h2593 : data <= 32'h67800000;
	16'h2594 : data <= 32'h130101fd;
	16'h2595 : data <= 32'h23261102;
	16'h2596 : data <= 32'h23248102;
	16'h2597 : data <= 32'h13040103;
	16'h2598 : data <= 32'h232ea4fc;
	16'h2599 : data <= 32'h8327c4fd;
	16'h259a : data <= 32'h03a70702;
	16'h259b : data <= 32'h93071000;
	16'h259c : data <= 32'h6316f70a;
	16'h259d : data <= 32'h8327c4fd;
	16'h259e : data <= 32'h83a7c700;
	16'h259f : data <= 32'h2326f4fe;
	16'h25a0 : data <= 32'h6f004004;
	16'h25a1 : data <= 32'h8327c4fd;
	16'h25a2 : data <= 32'h83a70700;
	16'h25a3 : data <= 32'h0327c4fd;
	16'h25a4 : data <= 32'h03274700;
	16'h25a5 : data <= 32'h03470700;
	16'h25a6 : data <= 32'h23a2e700;
	16'h25a7 : data <= 32'h8327c4fd;
	16'h25a8 : data <= 32'h83a74700;
	16'h25a9 : data <= 32'h13871700;
	16'h25aa : data <= 32'h8327c4fd;
	16'h25ab : data <= 32'h23a2e700;
	16'h25ac : data <= 32'h8327c4fd;
	16'h25ad : data <= 32'h83a7c700;
	16'h25ae : data <= 32'h1387f7ff;
	16'h25af : data <= 32'h8327c4fd;
	16'h25b0 : data <= 32'h23a6e700;
	16'h25b1 : data <= 32'h8327c4fd;
	16'h25b2 : data <= 32'h83a7c700;
	16'h25b3 : data <= 32'h638e0700;
	16'h25b4 : data <= 32'h8327c4fd;
	16'h25b5 : data <= 32'h83a70700;
	16'h25b6 : data <= 32'h83a7c700;
	16'h25b7 : data <= 32'h93d72700;
	16'h25b8 : data <= 32'h93f71700;
	16'h25b9 : data <= 32'he38007fa;
	16'h25ba : data <= 32'h8327c4fd;
	16'h25bb : data <= 32'h83a7c700;
	16'h25bc : data <= 32'h639a0702;
	16'h25bd : data <= 32'h8327c4fe;
	16'h25be : data <= 32'h63860702;
	16'h25bf : data <= 32'h8327c4fd;
	16'h25c0 : data <= 32'h83a74701;
	16'h25c1 : data <= 32'he7800700;
	16'h25c2 : data <= 32'h8327c4fd;
	16'h25c3 : data <= 32'h13072000;
	16'h25c4 : data <= 32'h23a0e702;
	16'h25c5 : data <= 32'h13000000;
	16'h25c6 : data <= 32'h6f00c000;
	16'h25c7 : data <= 32'h13000000;
	16'h25c8 : data <= 32'h6f008000;
	16'h25c9 : data <= 32'h13000000;
	16'h25ca : data <= 32'h8320c102;
	16'h25cb : data <= 32'h03248102;
	16'h25cc : data <= 32'h13010103;
	16'h25cd : data <= 32'h67800000;
	16'h25ce : data <= 32'h130101fd;
	16'h25cf : data <= 32'h23261102;
	16'h25d0 : data <= 32'h23248102;
	16'h25d1 : data <= 32'h13040103;
	16'h25d2 : data <= 32'h232ea4fc;
	16'h25d3 : data <= 32'h8327c4fd;
	16'h25d4 : data <= 32'h03a7c701;
	16'h25d5 : data <= 32'h93071000;
	16'h25d6 : data <= 32'h6318f70a;
	16'h25d7 : data <= 32'h8327c4fd;
	16'h25d8 : data <= 32'h83a70701;
	16'h25d9 : data <= 32'h2326f4fe;
	16'h25da : data <= 32'h6f008004;
	16'h25db : data <= 32'h8327c4fd;
	16'h25dc : data <= 32'h83a78700;
	16'h25dd : data <= 32'h0327c4fd;
	16'h25de : data <= 32'h03270700;
	16'h25df : data <= 32'h03278700;
	16'h25e0 : data <= 32'h1377f70f;
	16'h25e1 : data <= 32'h2380e700;
	16'h25e2 : data <= 32'h8327c4fd;
	16'h25e3 : data <= 32'h83a78700;
	16'h25e4 : data <= 32'h13871700;
	16'h25e5 : data <= 32'h8327c4fd;
	16'h25e6 : data <= 32'h23a4e700;
	16'h25e7 : data <= 32'h8327c4fd;
	16'h25e8 : data <= 32'h83a70701;
	16'h25e9 : data <= 32'h1387f7ff;
	16'h25ea : data <= 32'h8327c4fd;
	16'h25eb : data <= 32'h23a8e700;
	16'h25ec : data <= 32'h8327c4fd;
	16'h25ed : data <= 32'h83a70701;
	16'h25ee : data <= 32'h638e0700;
	16'h25ef : data <= 32'h8327c4fd;
	16'h25f0 : data <= 32'h83a70700;
	16'h25f1 : data <= 32'h83a7c700;
	16'h25f2 : data <= 32'h93d75700;
	16'h25f3 : data <= 32'h93f71700;
	16'h25f4 : data <= 32'he38e07f8;
	16'h25f5 : data <= 32'h8327c4fd;
	16'h25f6 : data <= 32'h83a70701;
	16'h25f7 : data <= 32'h639a0702;
	16'h25f8 : data <= 32'h8327c4fe;
	16'h25f9 : data <= 32'h63860702;
	16'h25fa : data <= 32'h8327c4fd;
	16'h25fb : data <= 32'h83a78701;
	16'h25fc : data <= 32'he7800700;
	16'h25fd : data <= 32'h8327c4fd;
	16'h25fe : data <= 32'h13072000;
	16'h25ff : data <= 32'h23aee700;
	16'h2600 : data <= 32'h13000000;
	16'h2601 : data <= 32'h6f00c000;
	16'h2602 : data <= 32'h13000000;
	16'h2603 : data <= 32'h6f008000;
	16'h2604 : data <= 32'h13000000;
	16'h2605 : data <= 32'h8320c102;
	16'h2606 : data <= 32'h03248102;
	16'h2607 : data <= 32'h13010103;
	16'h2608 : data <= 32'h67800000;
	16'h2609 : data <= 32'h4743433a;
	16'h260a : data <= 32'h2028474e;
	16'h260b : data <= 32'h55292035;
	16'h260c : data <= 32'h2e332e30;
	16'h260d : data <= 32'h00800080;
	16'h260e : data <= 32'h02000000;
	16'h260f : data <= 32'h02000000;
	16'h2610 : data <= 32'h00100080;
	16'h2611 : data <= 32'h03000000;
	16'h2612 : data <= 32'hFF;
	16'h3d : data <= 32'h4c990000;
	16'h2613 : data <= 32'h13000000;
	16'h2614 : data <= 32'h13000000;
	16'h2615 : data <= 32'h13000000;
	16'h2616 : data <= 32'h13000000;
	16'h2617 : data <= 32'h13000000;
	16'h2618 : data <= 32'h13000000;
	16'h2619 : data <= 32'h13000000;
	16'h261a : data <= 32'h13000000;
	16'h261b : data <= 32'h13000000;
	16'h261c : data <= 32'h13000000;
	16'h261d : data <= 32'h13000000;
	16'h261e : data <= 32'h13000000;
	16'h261f : data <= 32'h13000000;
	16'h2620 : data <= 32'h13000000;
	16'h2621 : data <= 32'h13000000;
	16'h2622 : data <= 32'h13000000;
	16'h2623 : data <= 32'h13000000;
	16'h2624 : data <= 32'h13000000;
	16'h2625 : data <= 32'h13000000;
	16'h2626 : data <= 32'h13000000;
	16'h2627 : data <= 32'h13000000;
	16'h2628 : data <= 32'h13000000;
	16'h2629 : data <= 32'h13000000;
	16'h262a : data <= 32'h13000000;
	16'h262b : data <= 32'h13000000;
	16'h262c : data <= 32'h13000000;
	16'h262d : data <= 32'h13000000;
	16'h262e : data <= 32'h13000000;
	16'h262f : data <= 32'h13000000;
	16'h2630 : data <= 32'h13000000;
	16'h2631 : data <= 32'h13000000;
	16'h2632 : data <= 32'h13000000;
	16'h2633 : data <= 32'h13000000;
	16'h2634 : data <= 32'h13000000;
	16'h2635 : data <= 32'h13000000;
	16'h2636 : data <= 32'h13000000;
	16'h2637 : data <= 32'h13000000;
	16'h2638 : data <= 32'h13000000;
	16'h2639 : data <= 32'h13000000;
	16'h263a : data <= 32'h13000000;
	16'h263b : data <= 32'h13000000;
	16'h263c : data <= 32'h13000000;
	16'h263d : data <= 32'h13000000;
	16'h263e : data <= 32'h13000000;
	16'h263f : data <= 32'h13000000;
	16'h2640 : data <= 32'h13000000;
	16'h2641 : data <= 32'h13000000;
	16'h2642 : data <= 32'h13000000;
	16'h2643 : data <= 32'h1301c1ff;
	16'h2644 : data <= 32'h23201100;
	16'h2645 : data <= 32'hef004006;
	16'h2646 : data <= 32'h83200100;
	16'h2647 : data <= 32'h13014100;
	16'h2648 : data <= 32'h73000010;
	16'h2649 : data <= 32'h13000000;
	16'h264a : data <= 32'h13000000;
	16'h264b : data <= 32'h13000000;
	16'h264c : data <= 32'h13000000;
	16'h264d : data <= 32'h13000000;
	16'h264e : data <= 32'h13000000;
	16'h264f : data <= 32'h13000000;
	16'h2650 : data <= 32'h13000000;
	16'h2651 : data <= 32'h13000000;
	16'h2652 : data <= 32'h13000000;
	16'h2653 : data <= 32'h13610000;
	16'h2654 : data <= 32'h1301c1ff;
	16'h2655 : data <= 32'h9362c000;
	16'h2656 : data <= 32'h9392c201;
	16'h2657 : data <= 32'h13630000;
	16'h2658 : data <= 32'h1303f3ff;
	16'h2659 : data <= 32'hb3c26200;
	16'h265a : data <= 32'h33715100;
	16'h265b : data <= 32'h97020000;
	16'h265c : data <= 32'h9382c27a;
	16'h265d : data <= 32'h67800200;
	16'h265e : data <= 32'h1301c1ff;
	16'h265f : data <= 32'h23201100;
	16'h2660 : data <= 32'h232ef1ff;
	16'h2661 : data <= 32'h232ce1ff;
	16'h2662 : data <= 32'h232ad1ff;
	16'h2663 : data <= 32'h2328c1ff;
	16'h2664 : data <= 32'h2326b1ff;
	16'h2665 : data <= 32'h2324a1ff;
	16'h2666 : data <= 32'h232291ff;
	16'h2667 : data <= 32'h232081ff;
	16'h2668 : data <= 32'h232e71fd;
	16'h2669 : data <= 32'h232c61fd;
	16'h266a : data <= 32'h232a51fd;
	16'h266b : data <= 32'h232841fd;
	16'h266c : data <= 32'h232631fd;
	16'h266d : data <= 32'h232421fd;
	16'h266e : data <= 32'h232211fd;
	16'h266f : data <= 32'h232001fd;
	16'h2670 : data <= 32'h232ef1fa;
	16'h2671 : data <= 32'h232ce1fa;
	16'h2672 : data <= 32'h232ad1fa;
	16'h2673 : data <= 32'h2328c1fa;
	16'h2674 : data <= 32'h2326b1fa;
	16'h2675 : data <= 32'h2324a1fa;
	16'h2676 : data <= 32'h232291fa;
	16'h2677 : data <= 32'h232081fa;
	16'h2678 : data <= 32'h232e71f8;
	16'h2679 : data <= 32'h232c61f8;
	16'h267a : data <= 32'h232a51f8;
	16'h267b : data <= 32'h232841f8;
	16'h267c : data <= 32'h232631f8;
	16'h267d : data <= 32'h232421f8;
	16'h267e : data <= 32'h232211f8;
	16'h267f : data <= 32'h232001f8;
	16'h2680 : data <= 32'h130101f8;
	16'h2681 : data <= 32'h93050100;
	16'h2682 : data <= 32'h73261034;
	16'h2683 : data <= 32'hf3263034;
	16'h2684 : data <= 32'h73252034;
	16'h2685 : data <= 32'h93020500;
	16'h2686 : data <= 32'h93d2f201;
	16'h2687 : data <= 32'h63860200;
	16'h2688 : data <= 32'hef004009;
	16'h2689 : data <= 32'h6f004001;
	16'h268a : data <= 32'hef00400d;
	16'h268b : data <= 32'hf3221034;
	16'h268c : data <= 32'h93824200;
	16'h268d : data <= 32'h73901234;
	16'h268e : data <= 32'h832fc107;
	16'h268f : data <= 32'h032f8107;
	16'h2690 : data <= 32'h832e4107;
	16'h2691 : data <= 32'h032e0107;
	16'h2692 : data <= 32'h832dc106;
	16'h2693 : data <= 32'h032d8106;
	16'h2694 : data <= 32'h832c4106;
	16'h2695 : data <= 32'h032c0106;
	16'h2696 : data <= 32'h832bc105;
	16'h2697 : data <= 32'h032b8105;
	16'h2698 : data <= 32'h832a4105;
	16'h2699 : data <= 32'h032a0105;
	16'h269a : data <= 32'h8329c104;
	16'h269b : data <= 32'h03298104;
	16'h269c : data <= 32'h83284104;
	16'h269d : data <= 32'h03280104;
	16'h269e : data <= 32'h8327c103;
	16'h269f : data <= 32'h03278103;
	16'h26a0 : data <= 32'h83264103;
	16'h26a1 : data <= 32'h03260103;
	16'h26a2 : data <= 32'h8325c102;
	16'h26a3 : data <= 32'h03258102;
	16'h26a4 : data <= 32'h83244102;
	16'h26a5 : data <= 32'h03240102;
	16'h26a6 : data <= 32'h8323c101;
	16'h26a7 : data <= 32'h03238101;
	16'h26a8 : data <= 32'h83224101;
	16'h26a9 : data <= 32'h13010108;
	16'h26aa : data <= 32'h83200100;
	16'h26ab : data <= 32'h13014100;
	16'h26ac : data <= 32'h67800000;
	16'h26ad : data <= 32'h130101fe;
	16'h26ae : data <= 32'h232e8100;
	16'h26af : data <= 32'h13040102;
	16'h26b0 : data <= 32'h2326a4fe;
	16'h26b1 : data <= 32'h13000000;
	16'h26b2 : data <= 32'h0324c101;
	16'h26b3 : data <= 32'h13010102;
	16'h26b4 : data <= 32'h67800000;
	16'h26b5 : data <= 32'h130101fe;
	16'h26b6 : data <= 32'h232e8100;
	16'h26b7 : data <= 32'h13040102;
	16'h26b8 : data <= 32'h2326a4fe;
	16'h26b9 : data <= 32'h8327c4fe;
	16'h26ba : data <= 32'hb307f040;
	16'h26bb : data <= 32'h13850700;
	16'h26bc : data <= 32'h0324c101;
	16'h26bd : data <= 32'h13010102;
	16'h26be : data <= 32'h67800000;
	16'h26bf : data <= 32'h130101fb;
	16'h26c0 : data <= 32'h23261104;
	16'h26c1 : data <= 32'h23248104;
	16'h26c2 : data <= 32'h23229104;
	16'h26c3 : data <= 32'h13040105;
	16'h26c4 : data <= 32'h232ea4fa;
	16'h26c5 : data <= 32'h232cb4fa;
	16'h26c6 : data <= 32'h232ac4fa;
	16'h26c7 : data <= 32'h2328d4fa;
	16'h26c8 : data <= 32'h0327c4fb;
	16'h26c9 : data <= 32'h93072000;
	16'h26ca : data <= 32'h6312f752;
	16'h26cb : data <= 32'h832744fb;
	16'h26cc : data <= 32'h83a70700;
	16'h26cd : data <= 32'h2326f4fe;
	16'h26ce : data <= 32'h8327c4fe;
	16'h26cf : data <= 32'h93f7f707;
	16'h26d0 : data <= 32'h2324f4fe;
	16'h26d1 : data <= 32'h0327c4fe;
	16'h26d2 : data <= 32'hb7170000;
	16'h26d3 : data <= 32'h938707f8;
	16'h26d4 : data <= 32'hb377f700;
	16'h26d5 : data <= 32'h93d77740;
	16'h26d6 : data <= 32'h2322f4fe;
	16'h26d7 : data <= 32'h0327c4fe;
	16'h26d8 : data <= 32'hb7870f00;
	16'h26d9 : data <= 32'hb377f700;
	16'h26da : data <= 32'h93d7f740;
	16'h26db : data <= 32'h2320f4fe;
	16'h26dc : data <= 32'h0327c4fe;
	16'h26dd : data <= 32'hb707f001;
	16'h26de : data <= 32'hb377f700;
	16'h26df : data <= 32'h93d74741;
	16'h26e0 : data <= 32'h232ef4fc;
	16'h26e1 : data <= 32'h0327c4fe;
	16'h26e2 : data <= 32'hb7770000;
	16'h26e3 : data <= 32'hb377f700;
	16'h26e4 : data <= 32'h93d7c740;
	16'h26e5 : data <= 32'h232cf4fc;
	16'h26e6 : data <= 32'h8327c4fe;
	16'h26e7 : data <= 32'h93d79701;
	16'h26e8 : data <= 32'h232af4fc;
	16'h26e9 : data <= 32'h032784fe;
	16'h26ea : data <= 32'h93073003;
	16'h26eb : data <= 32'h6310f74a;
	16'h26ec : data <= 32'h032744fd;
	16'h26ed : data <= 32'h93071000;
	16'h26ee : data <= 32'h631af748;
	16'h26ef : data <= 32'h832784fd;
	16'h26f0 : data <= 32'h63960704;
	16'h26f1 : data <= 32'h8327c4fd;
	16'h26f2 : data <= 32'h93972700;
	16'h26f3 : data <= 32'h032784fb;
	16'h26f4 : data <= 32'hb307f700;
	16'h26f5 : data <= 32'h83a60700;
	16'h26f6 : data <= 32'h832704fe;
	16'h26f7 : data <= 32'h93972700;
	16'h26f8 : data <= 32'h032784fb;
	16'h26f9 : data <= 32'hb307f700;
	16'h26fa : data <= 32'h83a50700;
	16'h26fb : data <= 32'h832744fe;
	16'h26fc : data <= 32'h93972700;
	16'h26fd : data <= 32'h032784fb;
	16'h26fe : data <= 32'hb307f700;
	16'h26ff : data <= 32'h13860700;
	16'h2700 : data <= 32'h13850600;
	16'h2701 : data <= 32'hef000046;
	16'h2702 : data <= 32'h6f004044;
	16'h2703 : data <= 32'h032784fd;
	16'h2704 : data <= 32'h93071000;
	16'h2705 : data <= 32'h630cf742;
	16'h2706 : data <= 32'h032784fd;
	16'h2707 : data <= 32'h93072000;
	16'h2708 : data <= 32'h6306f742;
	16'h2709 : data <= 32'h032784fd;
	16'h270a : data <= 32'h93073000;
	16'h270b : data <= 32'h6300f742;
	16'h270c : data <= 32'h032784fd;
	16'h270d : data <= 32'h93074000;
	16'h270e : data <= 32'h631cf716;
	16'h270f : data <= 32'h8327c4fd;
	16'h2710 : data <= 32'h93972700;
	16'h2711 : data <= 32'h032784fb;
	16'h2712 : data <= 32'hb307f700;
	16'h2713 : data <= 32'h83a70700;
	16'h2714 : data <= 32'h2328f4fc;
	16'h2715 : data <= 32'h832704fe;
	16'h2716 : data <= 32'h93972700;
	16'h2717 : data <= 32'h032784fb;
	16'h2718 : data <= 32'hb307f700;
	16'h2719 : data <= 32'h83a70700;
	16'h271a : data <= 32'h2326f4fc;
	16'h271b : data <= 32'h832704fd;
	16'h271c : data <= 32'h639c0700;
	16'h271d : data <= 32'h9307f0ff;
	16'h271e : data <= 32'h2324f4fc;
	16'h271f : data <= 32'h8327c4fc;
	16'h2720 : data <= 32'h2322f4fc;
	16'h2721 : data <= 32'h6f000011;
	16'h2722 : data <= 32'h0327c4fc;
	16'h2723 : data <= 32'hb7070080;
	16'h2724 : data <= 32'h6310f702;
	16'h2725 : data <= 32'h032704fd;
	16'h2726 : data <= 32'h9307f0ff;
	16'h2727 : data <= 32'h631af700;
	16'h2728 : data <= 32'h8327c4fc;
	16'h2729 : data <= 32'h2324f4fc;
	16'h272a : data <= 32'h232204fc;
	16'h272b : data <= 32'h6f00800e;
	16'h272c : data <= 32'h8327c4fc;
	16'h272d : data <= 32'h63d00704;
	16'h272e : data <= 32'h832704fd;
	16'h272f : data <= 32'h63dc0702;
	16'h2730 : data <= 32'h0325c4fc;
	16'h2731 : data <= 32'heff01fe1;
	16'h2732 : data <= 32'h93040500;
	16'h2733 : data <= 32'h032504fd;
	16'h2734 : data <= 32'heff05fe0;
	16'h2735 : data <= 32'h93050500;
	16'h2736 : data <= 32'h130744fc;
	16'h2737 : data <= 32'h930784fc;
	16'h2738 : data <= 32'h93060700;
	16'h2739 : data <= 32'h13860700;
	16'h273a : data <= 32'h13850400;
	16'h273b : data <= 32'hef00403c;
	16'h273c : data <= 32'h6f00400a;
	16'h273d : data <= 32'h8327c4fc;
	16'h273e : data <= 32'h63de0702;
	16'h273f : data <= 32'h0325c4fc;
	16'h2740 : data <= 32'heff05fdd;
	16'h2741 : data <= 32'h130744fc;
	16'h2742 : data <= 32'h930784fc;
	16'h2743 : data <= 32'h93060700;
	16'h2744 : data <= 32'h13860700;
	16'h2745 : data <= 32'h832504fd;
	16'h2746 : data <= 32'hef008039;
	16'h2747 : data <= 32'h832784fc;
	16'h2748 : data <= 32'h13850700;
	16'h2749 : data <= 32'heff01fdb;
	16'h274a : data <= 32'h93070500;
	16'h274b : data <= 32'h2324f4fc;
	16'h274c : data <= 32'h6f004006;
	16'h274d : data <= 32'h832704fd;
	16'h274e : data <= 32'h63d00704;
	16'h274f : data <= 32'h032504fd;
	16'h2750 : data <= 32'heff05fd9;
	16'h2751 : data <= 32'h93050500;
	16'h2752 : data <= 32'h130744fc;
	16'h2753 : data <= 32'h930784fc;
	16'h2754 : data <= 32'h93060700;
	16'h2755 : data <= 32'h13860700;
	16'h2756 : data <= 32'h0325c4fc;
	16'h2757 : data <= 32'hef004035;
	16'h2758 : data <= 32'h832784fc;
	16'h2759 : data <= 32'h13850700;
	16'h275a : data <= 32'heff0dfd6;
	16'h275b : data <= 32'h93070500;
	16'h275c : data <= 32'h2324f4fc;
	16'h275d : data <= 32'h6f000002;
	16'h275e : data <= 32'h130744fc;
	16'h275f : data <= 32'h930784fc;
	16'h2760 : data <= 32'h93060700;
	16'h2761 : data <= 32'h13860700;
	16'h2762 : data <= 32'h832504fd;
	16'h2763 : data <= 32'h0325c4fc;
	16'h2764 : data <= 32'hef000032;
	16'h2765 : data <= 32'h832744fe;
	16'h2766 : data <= 32'h93972700;
	16'h2767 : data <= 32'h032784fb;
	16'h2768 : data <= 32'hb307f700;
	16'h2769 : data <= 32'h032784fc;
	16'h276a : data <= 32'h23a0e700;
	16'h276b : data <= 32'h6f00002a;
	16'h276c : data <= 32'h032784fd;
	16'h276d : data <= 32'h93075000;
	16'h276e : data <= 32'h6314f708;
	16'h276f : data <= 32'h8327c4fd;
	16'h2770 : data <= 32'h93972700;
	16'h2771 : data <= 32'h032784fb;
	16'h2772 : data <= 32'hb307f700;
	16'h2773 : data <= 32'h83a70700;
	16'h2774 : data <= 32'h2328f4fc;
	16'h2775 : data <= 32'h832704fe;
	16'h2776 : data <= 32'h93972700;
	16'h2777 : data <= 32'h032784fb;
	16'h2778 : data <= 32'hb307f700;
	16'h2779 : data <= 32'h83a70700;
	16'h277a : data <= 32'h2326f4fc;
	16'h277b : data <= 32'h832704fd;
	16'h277c : data <= 32'h639c0700;
	16'h277d : data <= 32'h9307f0ff;
	16'h277e : data <= 32'h2324f4fc;
	16'h277f : data <= 32'h8327c4fc;
	16'h2780 : data <= 32'h2322f4fc;
	16'h2781 : data <= 32'h6f000002;
	16'h2782 : data <= 32'h130744fc;
	16'h2783 : data <= 32'h930784fc;
	16'h2784 : data <= 32'h93060700;
	16'h2785 : data <= 32'h13860700;
	16'h2786 : data <= 32'h832504fd;
	16'h2787 : data <= 32'h0325c4fc;
	16'h2788 : data <= 32'hef000029;
	16'h2789 : data <= 32'h832744fe;
	16'h278a : data <= 32'h93972700;
	16'h278b : data <= 32'h032784fb;
	16'h278c : data <= 32'hb307f700;
	16'h278d : data <= 32'h032784fc;
	16'h278e : data <= 32'h23a0e700;
	16'h278f : data <= 32'h6f000021;
	16'h2790 : data <= 32'h032784fd;
	16'h2791 : data <= 32'h93076000;
	16'h2792 : data <= 32'h631cf716;
	16'h2793 : data <= 32'h8327c4fd;
	16'h2794 : data <= 32'h93972700;
	16'h2795 : data <= 32'h032784fb;
	16'h2796 : data <= 32'hb307f700;
	16'h2797 : data <= 32'h83a70700;
	16'h2798 : data <= 32'h2328f4fc;
	16'h2799 : data <= 32'h832704fe;
	16'h279a : data <= 32'h93972700;
	16'h279b : data <= 32'h032784fb;
	16'h279c : data <= 32'hb307f700;
	16'h279d : data <= 32'h83a70700;
	16'h279e : data <= 32'h2326f4fc;
	16'h279f : data <= 32'h832704fd;
	16'h27a0 : data <= 32'h639c0700;
	16'h27a1 : data <= 32'h9307f0ff;
	16'h27a2 : data <= 32'h2324f4fc;
	16'h27a3 : data <= 32'h8327c4fc;
	16'h27a4 : data <= 32'h2322f4fc;
	16'h27a5 : data <= 32'h6f000011;
	16'h27a6 : data <= 32'h0327c4fc;
	16'h27a7 : data <= 32'hb7070080;
	16'h27a8 : data <= 32'h6310f702;
	16'h27a9 : data <= 32'h032704fd;
	16'h27aa : data <= 32'h9307f0ff;
	16'h27ab : data <= 32'h631af700;
	16'h27ac : data <= 32'h8327c4fc;
	16'h27ad : data <= 32'h2324f4fc;
	16'h27ae : data <= 32'h232204fc;
	16'h27af : data <= 32'h6f00800e;
	16'h27b0 : data <= 32'h8327c4fc;
	16'h27b1 : data <= 32'h63d00704;
	16'h27b2 : data <= 32'h832704fd;
	16'h27b3 : data <= 32'h63dc0702;
	16'h27b4 : data <= 32'h0325c4fc;
	16'h27b5 : data <= 32'heff01fc0;
	16'h27b6 : data <= 32'h93040500;
	16'h27b7 : data <= 32'h032504fd;
	16'h27b8 : data <= 32'heff05fbf;
	16'h27b9 : data <= 32'h93050500;
	16'h27ba : data <= 32'h130744fc;
	16'h27bb : data <= 32'h930784fc;
	16'h27bc : data <= 32'h93060700;
	16'h27bd : data <= 32'h13860700;
	16'h27be : data <= 32'h13850400;
	16'h27bf : data <= 32'hef00401b;
	16'h27c0 : data <= 32'h6f00400a;
	16'h27c1 : data <= 32'h8327c4fc;
	16'h27c2 : data <= 32'h63de0702;
	16'h27c3 : data <= 32'h0325c4fc;
	16'h27c4 : data <= 32'heff05fbc;
	16'h27c5 : data <= 32'h130744fc;
	16'h27c6 : data <= 32'h930784fc;
	16'h27c7 : data <= 32'h93060700;
	16'h27c8 : data <= 32'h13860700;
	16'h27c9 : data <= 32'h832504fd;
	16'h27ca : data <= 32'hef008018;
	16'h27cb : data <= 32'h832744fc;
	16'h27cc : data <= 32'h13850700;
	16'h27cd : data <= 32'heff01fba;
	16'h27ce : data <= 32'h93070500;
	16'h27cf : data <= 32'h2322f4fc;
	16'h27d0 : data <= 32'h6f004006;
	16'h27d1 : data <= 32'h832704fd;
	16'h27d2 : data <= 32'h63d00704;
	16'h27d3 : data <= 32'h032504fd;
	16'h27d4 : data <= 32'heff05fb8;
	16'h27d5 : data <= 32'h93050500;
	16'h27d6 : data <= 32'h130744fc;
	16'h27d7 : data <= 32'h930784fc;
	16'h27d8 : data <= 32'h93060700;
	16'h27d9 : data <= 32'h13860700;
	16'h27da : data <= 32'h0325c4fc;
	16'h27db : data <= 32'hef004014;
	16'h27dc : data <= 32'h832744fc;
	16'h27dd : data <= 32'h13850700;
	16'h27de : data <= 32'heff0dfb5;
	16'h27df : data <= 32'h93070500;
	16'h27e0 : data <= 32'h2322f4fc;
	16'h27e1 : data <= 32'h6f000002;
	16'h27e2 : data <= 32'h130744fc;
	16'h27e3 : data <= 32'h930784fc;
	16'h27e4 : data <= 32'h93060700;
	16'h27e5 : data <= 32'h13860700;
	16'h27e6 : data <= 32'h832504fd;
	16'h27e7 : data <= 32'h0325c4fc;
	16'h27e8 : data <= 32'hef000011;
	16'h27e9 : data <= 32'h832744fe;
	16'h27ea : data <= 32'h93972700;
	16'h27eb : data <= 32'h032784fb;
	16'h27ec : data <= 32'hb307f700;
	16'h27ed : data <= 32'h032744fc;
	16'h27ee : data <= 32'h23a0e700;
	16'h27ef : data <= 32'h6f000009;
	16'h27f0 : data <= 32'h032784fd;
	16'h27f1 : data <= 32'h93077000;
	16'h27f2 : data <= 32'h6312f708;
	16'h27f3 : data <= 32'h8327c4fd;
	16'h27f4 : data <= 32'h93972700;
	16'h27f5 : data <= 32'h032784fb;
	16'h27f6 : data <= 32'hb307f700;
	16'h27f7 : data <= 32'h83a70700;
	16'h27f8 : data <= 32'h2328f4fc;
	16'h27f9 : data <= 32'h832704fe;
	16'h27fa : data <= 32'h93972700;
	16'h27fb : data <= 32'h032784fb;
	16'h27fc : data <= 32'hb307f700;
	16'h27fd : data <= 32'h83a70700;
	16'h27fe : data <= 32'h2326f4fc;
	16'h27ff : data <= 32'h832704fd;
	16'h2800 : data <= 32'h639c0700;
	16'h2801 : data <= 32'h9307f0ff;
	16'h2802 : data <= 32'h2324f4fc;
	16'h2803 : data <= 32'h8327c4fc;
	16'h2804 : data <= 32'h2322f4fc;
	16'h2805 : data <= 32'h6f000002;
	16'h2806 : data <= 32'h130744fc;
	16'h2807 : data <= 32'h930784fc;
	16'h2808 : data <= 32'h93060700;
	16'h2809 : data <= 32'h13860700;
	16'h280a : data <= 32'h832504fd;
	16'h280b : data <= 32'h0325c4fc;
	16'h280c : data <= 32'hef000008;
	16'h280d : data <= 32'h832744fe;
	16'h280e : data <= 32'h93972700;
	16'h280f : data <= 32'h032784fb;
	16'h2810 : data <= 32'hb307f700;
	16'h2811 : data <= 32'h032744fc;
	16'h2812 : data <= 32'h23a0e700;
	16'h2813 : data <= 32'h13000000;
	16'h2814 : data <= 32'h8320c104;
	16'h2815 : data <= 32'h03248104;
	16'h2816 : data <= 32'h83244104;
	16'h2817 : data <= 32'h13010105;
	16'h2818 : data <= 32'h67800000;
	16'h2819 : data <= 32'h130101fe;
	16'h281a : data <= 32'h232e8100;
	16'h281b : data <= 32'h13040102;
	16'h281c : data <= 32'h2326a4fe;
	16'h281d : data <= 32'h2324b4fe;
	16'h281e : data <= 32'h2322c4fe;
	16'h281f : data <= 32'h93020500;
	16'h2820 : data <= 32'h13050000;
	16'h2821 : data <= 32'h13f31500;
	16'h2822 : data <= 32'h63040300;
	16'h2823 : data <= 32'h3385a200;
	16'h2824 : data <= 32'h93921200;
	16'h2825 : data <= 32'h93d51500;
	16'h2826 : data <= 32'he39605fe;
	16'h2827 : data <= 32'h2320a600;
	16'h2828 : data <= 32'h13000000;
	16'h2829 : data <= 32'h0324c101;
	16'h282a : data <= 32'h13010102;
	16'h282b : data <= 32'h67800000;
	16'h282c : data <= 32'h130101fe;
	16'h282d : data <= 32'h232e8100;
	16'h282e : data <= 32'h13040102;
	16'h282f : data <= 32'h2326a4fe;
	16'h2830 : data <= 32'h2324b4fe;
	16'h2831 : data <= 32'h2322c4fe;
	16'h2832 : data <= 32'h2320d4fe;
	16'h2833 : data <= 32'h93020000;
	16'h2834 : data <= 32'h13030000;
	16'h2835 : data <= 32'h130e1000;
	16'h2836 : data <= 32'h131efe01;
	16'h2837 : data <= 32'h13131300;
	16'h2838 : data <= 32'hb373c501;
	16'h2839 : data <= 32'h63840300;
	16'h283a : data <= 32'h13631300;
	16'h283b : data <= 32'h6346b300;
	16'h283c : data <= 32'h3303b340;
	16'h283d : data <= 32'hb3e2c201;
	16'h283e : data <= 32'h135e1e00;
	16'h283f : data <= 32'he3100efe;
	16'h2840 : data <= 32'h23205600;
	16'h2841 : data <= 32'h23a06600;
	16'h2842 : data <= 32'h13000000;
	16'h2843 : data <= 32'h0324c101;
	16'h2844 : data <= 32'h13010102;
	16'h2845 : data <= 32'h67800000;
	16'h2846 : data <= 32'h130101ff;
	16'h2847 : data <= 32'h23268100;
	16'h2848 : data <= 32'h13040101;
	16'h2849 : data <= 32'hb7070080;
	16'h284a : data <= 32'h23a40700;
	16'h284b : data <= 32'hb7070080;
	16'h284c : data <= 32'h37f7f0f0;
	16'h284d : data <= 32'h1307070f;
	16'h284e : data <= 32'h23a2e700;
	16'h284f : data <= 32'hb7b70000;
	16'h2850 : data <= 32'h93870768;
	16'h2851 : data <= 32'h13075005;
	16'h2852 : data <= 32'h23a0e700;
	16'h2853 : data <= 32'hb7c70000;
	16'h2854 : data <= 32'h93870788;
	16'h2855 : data <= 32'h13076006;
	16'h2856 : data <= 32'h23a0e700;
	16'h2857 : data <= 32'h93078002;
	16'h2858 : data <= 32'h23a00700;
	16'h2859 : data <= 32'hb7070080;
	16'h285a : data <= 32'h37f70000;
	16'h285b : data <= 32'h1307171f;
	16'h285c : data <= 32'h23a2e700;
	16'h285d : data <= 32'h93070002;
	16'h285e : data <= 32'h1307700c;
	16'h285f : data <= 32'h23a0e700;
	16'h2860 : data <= 32'hb7060080;
	16'h2861 : data <= 32'h93070002;
	16'h2862 : data <= 32'h03a70700;
	16'h2863 : data <= 32'h93070700;
	16'h2864 : data <= 32'h93978700;
	16'h2865 : data <= 32'hb387e700;
	16'h2866 : data <= 32'h13970701;
	16'h2867 : data <= 32'hb387e700;
	16'h2868 : data <= 32'h23a2f600;
	16'h2869 : data <= 32'h93074002;
	16'h286a : data <= 32'h13070002;
	16'h286b : data <= 32'h03270700;
	16'h286c : data <= 32'h13771700;
	16'h286d : data <= 32'h23a0e700;
	16'h286e : data <= 32'h93070002;
	16'h286f : data <= 32'h13070002;
	16'h2870 : data <= 32'h03270700;
	16'h2871 : data <= 32'h13571700;
	16'h2872 : data <= 32'h23a0e700;
	16'h2873 : data <= 32'h93074002;
	16'h2874 : data <= 32'h03a70700;
	16'h2875 : data <= 32'h93071000;
	16'h2876 : data <= 32'h631cf700;
	16'h2877 : data <= 32'h93070002;
	16'h2878 : data <= 32'h13070002;
	16'h2879 : data <= 32'h03270700;
	16'h287a : data <= 32'h1347870b;
	16'h287b : data <= 32'h23a0e700;
	16'h287c : data <= 32'h93078002;
	16'h287d : data <= 32'h23a00700;
	16'h287e : data <= 32'h13000000;
	16'h287f : data <= 32'h93078002;
	16'h2880 : data <= 32'h83a70700;
	16'h2881 : data <= 32'hb7060080;
	16'h2882 : data <= 32'h93070002;
	16'h2883 : data <= 32'h03a70700;
	16'h2884 : data <= 32'h93070700;
	16'h2885 : data <= 32'h93978700;
	16'h2886 : data <= 32'hb387e700;
	16'h2887 : data <= 32'h13970701;
	16'h2888 : data <= 32'hb387e700;
	16'h2889 : data <= 32'h23a2f600;
	16'h288a : data <= 32'h93070002;
	16'h288b : data <= 32'h03a70700;
	16'h288c : data <= 32'h9307f008;
	16'h288d : data <= 32'he318f7f6;
	16'h288e : data <= 32'hb7070080;
	16'h288f : data <= 32'h13074000;
	16'h2890 : data <= 32'h03270700;
	16'h2891 : data <= 32'h23a2e700;
	16'h2892 : data <= 32'h93078002;
	16'h2893 : data <= 32'h23a00700;
	16'h2894 : data <= 32'h6f004001;
	16'h2895 : data <= 32'h93078002;
	16'h2896 : data <= 32'h03a70700;
	16'h2897 : data <= 32'h13071700;
	16'h2898 : data <= 32'h23a0e700;
	16'h2899 : data <= 32'h93078002;
	16'h289a : data <= 32'h03a70700;
	16'h289b : data <= 32'hb7170000;
	16'h289c : data <= 32'h9387e7ff;
	16'h289d : data <= 32'he3f0e7fe;
	16'h289e : data <= 32'h93078002;
	16'h289f : data <= 32'h37070080;
	16'h28a0 : data <= 32'h03274700;
	16'h28a1 : data <= 32'h23a0e700;
	16'h28a2 : data <= 32'hb7070080;
	16'h28a3 : data <= 32'h13078002;
	16'h28a4 : data <= 32'h03270700;
	16'h28a5 : data <= 32'h23a2e700;
	16'h28a6 : data <= 32'h93070000;
	16'h28a7 : data <= 32'h83a70700;
	16'h28a8 : data <= 32'he38c07fc;
	16'h28a9 : data <= 32'h8322c000;
	16'h28aa : data <= 32'h67800200;
	16'h28ab : data <= 32'h13000000;
	16'h28ac : data <= 32'h13850700;
	16'h28ad : data <= 32'h0324c100;
	16'h28ae : data <= 32'h13010101;
	16'h28af : data <= 32'h67800000;
	16'h28b0 : data <= 32'h130101fd;
	16'h28b1 : data <= 32'h23268102;
	16'h28b2 : data <= 32'h13040103;
	16'h28b3 : data <= 32'h232ea4fc;
	16'h28b4 : data <= 32'h232cb4fc;
	16'h28b5 : data <= 32'h232ac4fc;
	16'h28b6 : data <= 32'h2328d4fc;
	16'h28b7 : data <= 32'h8327c4fd;
	16'h28b8 : data <= 32'h83a70700;
	16'h28b9 : data <= 32'h032784fd;
	16'h28ba : data <= 32'h23a4e700;
	16'h28bb : data <= 32'h8327c4fd;
	16'h28bc : data <= 32'h83a70700;
	16'h28bd : data <= 32'h032704fd;
	16'h28be : data <= 32'h23aae700;
	16'h28bf : data <= 32'h8327c4fd;
	16'h28c0 : data <= 32'h83a70700;
	16'h28c1 : data <= 32'h83a74700;
	16'h28c2 : data <= 32'h2326f4fe;
	16'h28c3 : data <= 32'h8327c4fe;
	16'h28c4 : data <= 32'h93f7e7ff;
	16'h28c5 : data <= 32'h2326f4fe;
	16'h28c6 : data <= 32'h8327c4fd;
	16'h28c7 : data <= 32'h83a70700;
	16'h28c8 : data <= 32'h032744fd;
	16'h28c9 : data <= 32'h93761700;
	16'h28ca : data <= 32'h0327c4fe;
	16'h28cb : data <= 32'h33e7e600;
	16'h28cc : data <= 32'h23a2e700;
	16'h28cd : data <= 32'h93070000;
	16'h28ce : data <= 32'h13850700;
	16'h28cf : data <= 32'h0324c102;
	16'h28d0 : data <= 32'h13010103;
	16'h28d1 : data <= 32'h67800000;
	16'h28d2 : data <= 32'h130101fc;
	16'h28d3 : data <= 32'h232e8102;
	16'h28d4 : data <= 32'h13040104;
	16'h28d5 : data <= 32'h2326a4fc;
	16'h28d6 : data <= 32'h2324b4fc;
	16'h28d7 : data <= 32'h2322c4fc;
	16'h28d8 : data <= 32'h232604fe;
	16'h28d9 : data <= 32'h032744fc;
	16'h28da : data <= 32'h93070004;
	16'h28db : data <= 32'h63f6e700;
	16'h28dc : data <= 32'h93070003;
	16'h28dd : data <= 32'h6f004020;
	16'h28de : data <= 32'h032744fc;
	16'h28df : data <= 32'h93070004;
	16'h28e0 : data <= 32'h631af702;
	16'h28e1 : data <= 32'h8327c4fc;
	16'h28e2 : data <= 32'h83a70700;
	16'h28e3 : data <= 32'h83a74700;
	16'h28e4 : data <= 32'h2322f4fe;
	16'h28e5 : data <= 32'h832744fe;
	16'h28e6 : data <= 32'h93f707fc;
	16'h28e7 : data <= 32'h2322f4fe;
	16'h28e8 : data <= 32'h8327c4fc;
	16'h28e9 : data <= 32'h83a70700;
	16'h28ea : data <= 32'h032744fe;
	16'h28eb : data <= 32'h23a2e700;
	16'h28ec : data <= 32'h6f000004;
	16'h28ed : data <= 32'h8327c4fc;
	16'h28ee : data <= 32'h83a70700;
	16'h28ef : data <= 32'h83a74700;
	16'h28f0 : data <= 32'h2320f4fe;
	16'h28f1 : data <= 32'h832704fe;
	16'h28f2 : data <= 32'h93f707fc;
	16'h28f3 : data <= 32'h2320f4fe;
	16'h28f4 : data <= 32'h8327c4fc;
	16'h28f5 : data <= 32'h83a70700;
	16'h28f6 : data <= 32'h032744fc;
	16'h28f7 : data <= 32'h13172700;
	16'h28f8 : data <= 32'h9376f70f;
	16'h28f9 : data <= 32'h032704fe;
	16'h28fa : data <= 32'h33e7e600;
	16'h28fb : data <= 32'h23a2e700;
	16'h28fc : data <= 32'h8327c4fc;
	16'h28fd : data <= 32'h83a70700;
	16'h28fe : data <= 32'h83a74700;
	16'h28ff : data <= 32'h232ef4fc;
	16'h2900 : data <= 32'h8327c4fd;
	16'h2901 : data <= 32'h93f7e7ff;
	16'h2902 : data <= 32'h232ef4fc;
	16'h2903 : data <= 32'h8327c4fc;
	16'h2904 : data <= 32'h83a70700;
	16'h2905 : data <= 32'h0327c4fd;
	16'h2906 : data <= 32'h13670710;
	16'h2907 : data <= 32'h23a2e700;
	16'h2908 : data <= 32'h8327c4fc;
	16'h2909 : data <= 32'h83a70700;
	16'h290a : data <= 32'h83a74700;
	16'h290b : data <= 32'h232cf4fc;
	16'h290c : data <= 32'h832784fd;
	16'h290d : data <= 32'h93f7e7ff;
	16'h290e : data <= 32'h232cf4fc;
	16'h290f : data <= 32'h8327c4fc;
	16'h2910 : data <= 32'h83a70700;
	16'h2911 : data <= 32'h032784fd;
	16'h2912 : data <= 32'h23a2e700;
	16'h2913 : data <= 32'h6f008002;
	16'h2914 : data <= 32'h8327c4fc;
	16'h2915 : data <= 32'h03a70700;
	16'h2916 : data <= 32'h8327c4fe;
	16'h2917 : data <= 32'h93861700;
	16'h2918 : data <= 32'h2326d4fe;
	16'h2919 : data <= 32'h832684fc;
	16'h291a : data <= 32'hb387f600;
	16'h291b : data <= 32'h83c70700;
	16'h291c : data <= 32'h2320f700;
	16'h291d : data <= 32'h0327c4fe;
	16'h291e : data <= 32'h832744fc;
	16'h291f : data <= 32'h637ef700;
	16'h2920 : data <= 32'h8327c4fc;
	16'h2921 : data <= 32'h83a70700;
	16'h2922 : data <= 32'h83a70701;
	16'h2923 : data <= 32'h93d7b700;
	16'h2924 : data <= 32'h93f71700;
	16'h2925 : data <= 32'he38e07fa;
	16'h2926 : data <= 32'h8327c4fc;
	16'h2927 : data <= 32'h83a70700;
	16'h2928 : data <= 32'h83a74700;
	16'h2929 : data <= 32'h232af4fc;
	16'h292a : data <= 32'h832744fd;
	16'h292b : data <= 32'h93f7e7ff;
	16'h292c : data <= 32'h232af4fc;
	16'h292d : data <= 32'h8327c4fc;
	16'h292e : data <= 32'h83a70700;
	16'h292f : data <= 32'h032744fd;
	16'h2930 : data <= 32'h13670720;
	16'h2931 : data <= 32'h23a2e700;
	16'h2932 : data <= 32'h8327c4fc;
	16'h2933 : data <= 32'h83a70700;
	16'h2934 : data <= 32'h83a70701;
	16'h2935 : data <= 32'h2324f4fe;
	16'h2936 : data <= 32'h6f000008;
	16'h2937 : data <= 32'h832784fe;
	16'h2938 : data <= 32'h93f71700;
	16'h2939 : data <= 32'h63860700;
	16'h293a : data <= 32'h93071003;
	16'h293b : data <= 32'h6f00c008;
	16'h293c : data <= 32'h832784fe;
	16'h293d : data <= 32'h93d73700;
	16'h293e : data <= 32'h93f71700;
	16'h293f : data <= 32'h63860700;
	16'h2940 : data <= 32'h93072003;
	16'h2941 : data <= 32'h6f004007;
	16'h2942 : data <= 32'h832784fe;
	16'h2943 : data <= 32'h93d7b700;
	16'h2944 : data <= 32'h93f71700;
	16'h2945 : data <= 32'h639a0702;
	16'h2946 : data <= 32'h0327c4fe;
	16'h2947 : data <= 32'h832744fc;
	16'h2948 : data <= 32'h6374f702;
	16'h2949 : data <= 32'h8327c4fc;
	16'h294a : data <= 32'h03a70700;
	16'h294b : data <= 32'h8327c4fe;
	16'h294c : data <= 32'h93861700;
	16'h294d : data <= 32'h2326d4fe;
	16'h294e : data <= 32'h832684fc;
	16'h294f : data <= 32'hb387f600;
	16'h2950 : data <= 32'h83c70700;
	16'h2951 : data <= 32'h2320f700;
	16'h2952 : data <= 32'h8327c4fc;
	16'h2953 : data <= 32'h83a70700;
	16'h2954 : data <= 32'h83a70701;
	16'h2955 : data <= 32'h2324f4fe;
	16'h2956 : data <= 32'h0327c4fe;
	16'h2957 : data <= 32'h832744fc;
	16'h2958 : data <= 32'he36ef7f6;
	16'h2959 : data <= 32'h832784fe;
	16'h295a : data <= 32'h93d72700;
	16'h295b : data <= 32'h93f71700;
	16'h295c : data <= 32'he38607f6;
	16'h295d : data <= 32'h93070000;
	16'h295e : data <= 32'h13850700;
	16'h295f : data <= 32'h0324c103;
	16'h2960 : data <= 32'h13010104;
	16'h2961 : data <= 32'h67800000;
	16'h2962 : data <= 32'h130101fc;
	16'h2963 : data <= 32'h232e8102;
	16'h2964 : data <= 32'h13040104;
	16'h2965 : data <= 32'h2326a4fc;
	16'h2966 : data <= 32'h2324b4fc;
	16'h2967 : data <= 32'h2322c4fc;
	16'h2968 : data <= 32'h232604fe;
	16'h2969 : data <= 32'h032744fc;
	16'h296a : data <= 32'h93070004;
	16'h296b : data <= 32'h63f6e700;
	16'h296c : data <= 32'h93070003;
	16'h296d : data <= 32'h6f00401e;
	16'h296e : data <= 32'h032744fc;
	16'h296f : data <= 32'h93070004;
	16'h2970 : data <= 32'h631af702;
	16'h2971 : data <= 32'h8327c4fc;
	16'h2972 : data <= 32'h83a70700;
	16'h2973 : data <= 32'h83a74700;
	16'h2974 : data <= 32'h2322f4fe;
	16'h2975 : data <= 32'h832744fe;
	16'h2976 : data <= 32'h93f707fc;
	16'h2977 : data <= 32'h2322f4fe;
	16'h2978 : data <= 32'h8327c4fc;
	16'h2979 : data <= 32'h83a70700;
	16'h297a : data <= 32'h032744fe;
	16'h297b : data <= 32'h23a2e700;
	16'h297c : data <= 32'h6f000004;
	16'h297d : data <= 32'h8327c4fc;
	16'h297e : data <= 32'h83a70700;
	16'h297f : data <= 32'h83a74700;
	16'h2980 : data <= 32'h2320f4fe;
	16'h2981 : data <= 32'h832704fe;
	16'h2982 : data <= 32'h93f707fc;
	16'h2983 : data <= 32'h2320f4fe;
	16'h2984 : data <= 32'h8327c4fc;
	16'h2985 : data <= 32'h83a70700;
	16'h2986 : data <= 32'h032744fc;
	16'h2987 : data <= 32'h13172700;
	16'h2988 : data <= 32'h9376f70f;
	16'h2989 : data <= 32'h032704fe;
	16'h298a : data <= 32'h33e7e600;
	16'h298b : data <= 32'h23a2e700;
	16'h298c : data <= 32'h8327c4fc;
	16'h298d : data <= 32'h83a70700;
	16'h298e : data <= 32'h83a74700;
	16'h298f : data <= 32'h232ef4fc;
	16'h2990 : data <= 32'h8327c4fd;
	16'h2991 : data <= 32'h93f7e7ff;
	16'h2992 : data <= 32'h232ef4fc;
	16'h2993 : data <= 32'h8327c4fc;
	16'h2994 : data <= 32'h83a70700;
	16'h2995 : data <= 32'h0327c4fd;
	16'h2996 : data <= 32'h23a2e700;
	16'h2997 : data <= 32'h8327c4fc;
	16'h2998 : data <= 32'h83a70700;
	16'h2999 : data <= 32'h83a74700;
	16'h299a : data <= 32'h232cf4fc;
	16'h299b : data <= 32'h832784fd;
	16'h299c : data <= 32'h93f7e7ff;
	16'h299d : data <= 32'h232cf4fc;
	16'h299e : data <= 32'h8327c4fc;
	16'h299f : data <= 32'h83a70700;
	16'h29a0 : data <= 32'h032784fd;
	16'h29a1 : data <= 32'h23a2e700;
	16'h29a2 : data <= 32'h6f004001;
	16'h29a3 : data <= 32'h8327c4fc;
	16'h29a4 : data <= 32'h83a70700;
	16'h29a5 : data <= 32'h83a7c700;
	16'h29a6 : data <= 32'h232af4fc;
	16'h29a7 : data <= 32'h8327c4fc;
	16'h29a8 : data <= 32'h83a70700;
	16'h29a9 : data <= 32'h83a70701;
	16'h29aa : data <= 32'h93d77700;
	16'h29ab : data <= 32'h93f71700;
	16'h29ac : data <= 32'he38e07fc;
	16'h29ad : data <= 32'h8327c4fc;
	16'h29ae : data <= 32'h83a70700;
	16'h29af : data <= 32'h83a74700;
	16'h29b0 : data <= 32'h2328f4fc;
	16'h29b1 : data <= 32'h832704fd;
	16'h29b2 : data <= 32'h93f7e7ff;
	16'h29b3 : data <= 32'h2328f4fc;
	16'h29b4 : data <= 32'h8327c4fc;
	16'h29b5 : data <= 32'h83a70700;
	16'h29b6 : data <= 32'h032704fd;
	16'h29b7 : data <= 32'h13670720;
	16'h29b8 : data <= 32'h23a2e700;
	16'h29b9 : data <= 32'h8327c4fc;
	16'h29ba : data <= 32'h83a70700;
	16'h29bb : data <= 32'h83a70701;
	16'h29bc : data <= 32'h2324f4fe;
	16'h29bd : data <= 32'h6f004008;
	16'h29be : data <= 32'h832784fe;
	16'h29bf : data <= 32'h93f71700;
	16'h29c0 : data <= 32'h63860700;
	16'h29c1 : data <= 32'h93071003;
	16'h29c2 : data <= 32'h6f000009;
	16'h29c3 : data <= 32'h832784fe;
	16'h29c4 : data <= 32'h93d73700;
	16'h29c5 : data <= 32'h93f71700;
	16'h29c6 : data <= 32'h63860700;
	16'h29c7 : data <= 32'h93072003;
	16'h29c8 : data <= 32'h6f008007;
	16'h29c9 : data <= 32'h832784fe;
	16'h29ca : data <= 32'h93d77700;
	16'h29cb : data <= 32'h93f71700;
	16'h29cc : data <= 32'h639c0702;
	16'h29cd : data <= 32'h0327c4fe;
	16'h29ce : data <= 32'h832744fc;
	16'h29cf : data <= 32'h6376f702;
	16'h29d0 : data <= 32'h8327c4fe;
	16'h29d1 : data <= 32'h13871700;
	16'h29d2 : data <= 32'h2326e4fe;
	16'h29d3 : data <= 32'h032784fc;
	16'h29d4 : data <= 32'hb307f700;
	16'h29d5 : data <= 32'h0327c4fc;
	16'h29d6 : data <= 32'h03270700;
	16'h29d7 : data <= 32'h0327c700;
	16'h29d8 : data <= 32'h1377f70f;
	16'h29d9 : data <= 32'h2380e700;
	16'h29da : data <= 32'h8327c4fc;
	16'h29db : data <= 32'h83a70700;
	16'h29dc : data <= 32'h83a70701;
	16'h29dd : data <= 32'h2324f4fe;
	16'h29de : data <= 32'h0327c4fe;
	16'h29df : data <= 32'h832744fc;
	16'h29e0 : data <= 32'he36cf7f6;
	16'h29e1 : data <= 32'h832784fe;
	16'h29e2 : data <= 32'h93d72700;
	16'h29e3 : data <= 32'h93f71700;
	16'h29e4 : data <= 32'he38407f6;
	16'h29e5 : data <= 32'h93070000;
	16'h29e6 : data <= 32'h13850700;
	16'h29e7 : data <= 32'h0324c103;
	16'h29e8 : data <= 32'h13010104;
	16'h29e9 : data <= 32'h67800000;
	16'h29ea : data <= 32'h130101fc;
	16'h29eb : data <= 32'h232e8102;
	16'h29ec : data <= 32'h13040104;
	16'h29ed : data <= 32'h2326a4fc;
	16'h29ee : data <= 32'h2324b4fc;
	16'h29ef : data <= 32'h2322c4fc;
	16'h29f0 : data <= 32'h2320d4fc;
	16'h29f1 : data <= 32'h232604fe;
	16'h29f2 : data <= 32'h032744fc;
	16'h29f3 : data <= 32'h93070004;
	16'h29f4 : data <= 32'h63f6e700;
	16'h29f5 : data <= 32'h93070003;
	16'h29f6 : data <= 32'h6f00801d;
	16'h29f7 : data <= 32'h032744fc;
	16'h29f8 : data <= 32'h93070004;
	16'h29f9 : data <= 32'h631af702;
	16'h29fa : data <= 32'h8327c4fc;
	16'h29fb : data <= 32'h83a70700;
	16'h29fc : data <= 32'h83a74700;
	16'h29fd : data <= 32'h2324f4fe;
	16'h29fe : data <= 32'h832784fe;
	16'h29ff : data <= 32'h93f707fc;
	16'h2a00 : data <= 32'h2324f4fe;
	16'h2a01 : data <= 32'h8327c4fc;
	16'h2a02 : data <= 32'h83a70700;
	16'h2a03 : data <= 32'h032784fe;
	16'h2a04 : data <= 32'h23a2e700;
	16'h2a05 : data <= 32'h6f000004;
	16'h2a06 : data <= 32'h8327c4fc;
	16'h2a07 : data <= 32'h83a70700;
	16'h2a08 : data <= 32'h83a74700;
	16'h2a09 : data <= 32'h2322f4fe;
	16'h2a0a : data <= 32'h832744fe;
	16'h2a0b : data <= 32'h93f707fc;
	16'h2a0c : data <= 32'h2322f4fe;
	16'h2a0d : data <= 32'h8327c4fc;
	16'h2a0e : data <= 32'h83a70700;
	16'h2a0f : data <= 32'h032744fc;
	16'h2a10 : data <= 32'h13172700;
	16'h2a11 : data <= 32'h9376f70f;
	16'h2a12 : data <= 32'h032744fe;
	16'h2a13 : data <= 32'h33e7e600;
	16'h2a14 : data <= 32'h23a2e700;
	16'h2a15 : data <= 32'h8327c4fc;
	16'h2a16 : data <= 32'h83a70700;
	16'h2a17 : data <= 32'h83a74700;
	16'h2a18 : data <= 32'h2320f4fe;
	16'h2a19 : data <= 32'h832704fe;
	16'h2a1a : data <= 32'h93f7e7ff;
	16'h2a1b : data <= 32'h2320f4fe;
	16'h2a1c : data <= 32'h8327c4fc;
	16'h2a1d : data <= 32'h83a70700;
	16'h2a1e : data <= 32'h032704fe;
	16'h2a1f : data <= 32'h13670710;
	16'h2a20 : data <= 32'h23a2e700;
	16'h2a21 : data <= 32'h8327c4fc;
	16'h2a22 : data <= 32'h83a70700;
	16'h2a23 : data <= 32'h83a74700;
	16'h2a24 : data <= 32'h232ef4fc;
	16'h2a25 : data <= 32'h8327c4fd;
	16'h2a26 : data <= 32'h93f7e7ff;
	16'h2a27 : data <= 32'h232ef4fc;
	16'h2a28 : data <= 32'h8327c4fc;
	16'h2a29 : data <= 32'h83a70700;
	16'h2a2a : data <= 32'h0327c4fd;
	16'h2a2b : data <= 32'h23a2e700;
	16'h2a2c : data <= 32'h6f000003;
	16'h2a2d : data <= 32'h8327c4fc;
	16'h2a2e : data <= 32'h83a70700;
	16'h2a2f : data <= 32'h032784fc;
	16'h2a30 : data <= 32'h03470700;
	16'h2a31 : data <= 32'h23a0e700;
	16'h2a32 : data <= 32'h832784fc;
	16'h2a33 : data <= 32'h93871700;
	16'h2a34 : data <= 32'h2324f4fc;
	16'h2a35 : data <= 32'h832744fc;
	16'h2a36 : data <= 32'h9387f7ff;
	16'h2a37 : data <= 32'h2322f4fc;
	16'h2a38 : data <= 32'h832744fc;
	16'h2a39 : data <= 32'h638e0700;
	16'h2a3a : data <= 32'h8327c4fc;
	16'h2a3b : data <= 32'h83a70700;
	16'h2a3c : data <= 32'h83a70701;
	16'h2a3d : data <= 32'h93d7b700;
	16'h2a3e : data <= 32'h93f71700;
	16'h2a3f : data <= 32'he38c07fa;
	16'h2a40 : data <= 32'h8327c4fc;
	16'h2a41 : data <= 32'h032784fc;
	16'h2a42 : data <= 32'h23a2e700;
	16'h2a43 : data <= 32'h8327c4fc;
	16'h2a44 : data <= 32'h032744fc;
	16'h2a45 : data <= 32'h23a4e700;
	16'h2a46 : data <= 32'h8327c4fc;
	16'h2a47 : data <= 32'h032704fc;
	16'h2a48 : data <= 32'h23a6e700;
	16'h2a49 : data <= 32'h6f008002;
	16'h2a4a : data <= 32'h8327c4fc;
	16'h2a4b : data <= 32'h03a70700;
	16'h2a4c : data <= 32'h8327c4fe;
	16'h2a4d : data <= 32'h93861700;
	16'h2a4e : data <= 32'h2326d4fe;
	16'h2a4f : data <= 32'h832684fc;
	16'h2a50 : data <= 32'hb387f600;
	16'h2a51 : data <= 32'h83c70700;
	16'h2a52 : data <= 32'h2320f700;
	16'h2a53 : data <= 32'h0327c4fe;
	16'h2a54 : data <= 32'h832744fc;
	16'h2a55 : data <= 32'h637ef700;
	16'h2a56 : data <= 32'h8327c4fc;
	16'h2a57 : data <= 32'h83a70700;
	16'h2a58 : data <= 32'h83a70701;
	16'h2a59 : data <= 32'h93d7b700;
	16'h2a5a : data <= 32'h93f71700;
	16'h2a5b : data <= 32'he38e07fa;
	16'h2a5c : data <= 32'h8327c4fc;
	16'h2a5d : data <= 32'h83a70700;
	16'h2a5e : data <= 32'h83a74700;
	16'h2a5f : data <= 32'h232cf4fc;
	16'h2a60 : data <= 32'h832784fd;
	16'h2a61 : data <= 32'h93f7e7ff;
	16'h2a62 : data <= 32'h232cf4fc;
	16'h2a63 : data <= 32'h8327c4fc;
	16'h2a64 : data <= 32'h83a70700;
	16'h2a65 : data <= 32'h032784fd;
	16'h2a66 : data <= 32'h13670720;
	16'h2a67 : data <= 32'h23a2e700;
	16'h2a68 : data <= 32'h8327c4fc;
	16'h2a69 : data <= 32'h13071000;
	16'h2a6a : data <= 32'h23a8e700;
	16'h2a6b : data <= 32'h93070000;
	16'h2a6c : data <= 32'h13850700;
	16'h2a6d : data <= 32'h0324c103;
	16'h2a6e : data <= 32'h13010104;
	16'h2a6f : data <= 32'h67800000;
	16'h2a70 : data <= 32'h130101fd;
	16'h2a71 : data <= 32'h23268102;
	16'h2a72 : data <= 32'h13040103;
	16'h2a73 : data <= 32'h232ea4fc;
	16'h2a74 : data <= 32'h232cb4fc;
	16'h2a75 : data <= 32'h232ac4fc;
	16'h2a76 : data <= 32'h232604fe;
	16'h2a77 : data <= 32'h8327c4fd;
	16'h2a78 : data <= 32'h83a70700;
	16'h2a79 : data <= 32'h83a74700;
	16'h2a7a : data <= 32'h2322f4fe;
	16'h2a7b : data <= 32'h832744fe;
	16'h2a7c : data <= 32'h93f7e7ff;
	16'h2a7d : data <= 32'h2322f4fe;
	16'h2a7e : data <= 32'h8327c4fd;
	16'h2a7f : data <= 32'h83a70700;
	16'h2a80 : data <= 32'h032744fe;
	16'h2a81 : data <= 32'h13672700;
	16'h2a82 : data <= 32'h23a2e700;
	16'h2a83 : data <= 32'h6f008002;
	16'h2a84 : data <= 32'h8327c4fd;
	16'h2a85 : data <= 32'h03a70700;
	16'h2a86 : data <= 32'h8327c4fe;
	16'h2a87 : data <= 32'h93861700;
	16'h2a88 : data <= 32'h2326d4fe;
	16'h2a89 : data <= 32'h832684fd;
	16'h2a8a : data <= 32'hb387f600;
	16'h2a8b : data <= 32'h83c70700;
	16'h2a8c : data <= 32'h2320f700;
	16'h2a8d : data <= 32'h0327c4fe;
	16'h2a8e : data <= 32'h832744fd;
	16'h2a8f : data <= 32'h637ef700;
	16'h2a90 : data <= 32'h8327c4fd;
	16'h2a91 : data <= 32'h83a70700;
	16'h2a92 : data <= 32'h83a70701;
	16'h2a93 : data <= 32'h93d7b700;
	16'h2a94 : data <= 32'h93f71700;
	16'h2a95 : data <= 32'he38e07fa;
	16'h2a96 : data <= 32'h8327c4fd;
	16'h2a97 : data <= 32'h83a70700;
	16'h2a98 : data <= 32'h83a70701;
	16'h2a99 : data <= 32'h2324f4fe;
	16'h2a9a : data <= 32'h6f008006;
	16'h2a9b : data <= 32'h832784fe;
	16'h2a9c : data <= 32'h93f71700;
	16'h2a9d : data <= 32'h63860700;
	16'h2a9e : data <= 32'h93071003;
	16'h2a9f : data <= 32'h6f004007;
	16'h2aa0 : data <= 32'h832784fe;
	16'h2aa1 : data <= 32'h93d7b700;
	16'h2aa2 : data <= 32'h93f71700;
	16'h2aa3 : data <= 32'h639a0702;
	16'h2aa4 : data <= 32'h0327c4fe;
	16'h2aa5 : data <= 32'h832744fd;
	16'h2aa6 : data <= 32'h6374f702;
	16'h2aa7 : data <= 32'h8327c4fd;
	16'h2aa8 : data <= 32'h03a70700;
	16'h2aa9 : data <= 32'h8327c4fe;
	16'h2aaa : data <= 32'h93861700;
	16'h2aab : data <= 32'h2326d4fe;
	16'h2aac : data <= 32'h832684fd;
	16'h2aad : data <= 32'hb387f600;
	16'h2aae : data <= 32'h83c70700;
	16'h2aaf : data <= 32'h2320f700;
	16'h2ab0 : data <= 32'h8327c4fd;
	16'h2ab1 : data <= 32'h83a70700;
	16'h2ab2 : data <= 32'h83a70701;
	16'h2ab3 : data <= 32'h2324f4fe;
	16'h2ab4 : data <= 32'h0327c4fe;
	16'h2ab5 : data <= 32'h832744fd;
	16'h2ab6 : data <= 32'he36af7f8;
	16'h2ab7 : data <= 32'h832784fe;
	16'h2ab8 : data <= 32'h93d72700;
	16'h2ab9 : data <= 32'h93f71700;
	16'h2aba : data <= 32'he38207f8;
	16'h2abb : data <= 32'h93070000;
	16'h2abc : data <= 32'h13850700;
	16'h2abd : data <= 32'h0324c102;
	16'h2abe : data <= 32'h13010103;
	16'h2abf : data <= 32'h67800000;
	16'h2ac0 : data <= 32'h130101fd;
	16'h2ac1 : data <= 32'h23268102;
	16'h2ac2 : data <= 32'h13040103;
	16'h2ac3 : data <= 32'h232ea4fc;
	16'h2ac4 : data <= 32'h232cb4fc;
	16'h2ac5 : data <= 32'h232ac4fc;
	16'h2ac6 : data <= 32'h232604fe;
	16'h2ac7 : data <= 32'h8327c4fd;
	16'h2ac8 : data <= 32'h83a70700;
	16'h2ac9 : data <= 32'h83a74700;
	16'h2aca : data <= 32'h2322f4fe;
	16'h2acb : data <= 32'h832744fe;
	16'h2acc : data <= 32'h93f7e7ff;
	16'h2acd : data <= 32'h2322f4fe;
	16'h2ace : data <= 32'h8327c4fd;
	16'h2acf : data <= 32'h83a70700;
	16'h2ad0 : data <= 32'h032744fe;
	16'h2ad1 : data <= 32'h13672700;
	16'h2ad2 : data <= 32'h23a2e700;
	16'h2ad3 : data <= 32'h6f004001;
	16'h2ad4 : data <= 32'h8327c4fd;
	16'h2ad5 : data <= 32'h83a70700;
	16'h2ad6 : data <= 32'h83a7c700;
	16'h2ad7 : data <= 32'h2320f4fe;
	16'h2ad8 : data <= 32'h8327c4fd;
	16'h2ad9 : data <= 32'h83a70700;
	16'h2ada : data <= 32'h83a70701;
	16'h2adb : data <= 32'h93d77700;
	16'h2adc : data <= 32'h93f71700;
	16'h2add : data <= 32'he38e07fc;
	16'h2ade : data <= 32'h8327c4fd;
	16'h2adf : data <= 32'h83a70700;
	16'h2ae0 : data <= 32'h83a70701;
	16'h2ae1 : data <= 32'h2324f4fe;
	16'h2ae2 : data <= 32'h6f00c006;
	16'h2ae3 : data <= 32'h832784fe;
	16'h2ae4 : data <= 32'h93f71700;
	16'h2ae5 : data <= 32'h63860700;
	16'h2ae6 : data <= 32'h93071003;
	16'h2ae7 : data <= 32'h6f008007;
	16'h2ae8 : data <= 32'h832784fe;
	16'h2ae9 : data <= 32'h93d77700;
	16'h2aea : data <= 32'h93f71700;
	16'h2aeb : data <= 32'h639c0702;
	16'h2aec : data <= 32'h0327c4fe;
	16'h2aed : data <= 32'h832744fd;
	16'h2aee : data <= 32'h6376f702;
	16'h2aef : data <= 32'h8327c4fe;
	16'h2af0 : data <= 32'h13871700;
	16'h2af1 : data <= 32'h2326e4fe;
	16'h2af2 : data <= 32'h032784fd;
	16'h2af3 : data <= 32'hb307f700;
	16'h2af4 : data <= 32'h0327c4fd;
	16'h2af5 : data <= 32'h03270700;
	16'h2af6 : data <= 32'h0327c700;
	16'h2af7 : data <= 32'h1377f70f;
	16'h2af8 : data <= 32'h2380e700;
	16'h2af9 : data <= 32'h8327c4fd;
	16'h2afa : data <= 32'h83a70700;
	16'h2afb : data <= 32'h83a70701;
	16'h2afc : data <= 32'h2324f4fe;
	16'h2afd : data <= 32'h0327c4fe;
	16'h2afe : data <= 32'h832744fd;
	16'h2aff : data <= 32'he368f7f8;
	16'h2b00 : data <= 32'h832784fe;
	16'h2b01 : data <= 32'h93d72700;
	16'h2b02 : data <= 32'h93f71700;
	16'h2b03 : data <= 32'he38007f8;
	16'h2b04 : data <= 32'h93070000;
	16'h2b05 : data <= 32'h13850700;
	16'h2b06 : data <= 32'h0324c102;
	16'h2b07 : data <= 32'h13010103;
	16'h2b08 : data <= 32'h67800000;
	16'h2b09 : data <= 32'h130101fd;
	16'h2b0a : data <= 32'h23268102;
	16'h2b0b : data <= 32'h13040103;
	16'h2b0c : data <= 32'h232ea4fc;
	16'h2b0d : data <= 32'h232cb4fc;
	16'h2b0e : data <= 32'h232ac4fc;
	16'h2b0f : data <= 32'h2328d4fc;
	16'h2b10 : data <= 32'h232604fe;
	16'h2b11 : data <= 32'h8327c4fd;
	16'h2b12 : data <= 32'h83a70700;
	16'h2b13 : data <= 32'h83a74700;
	16'h2b14 : data <= 32'h2324f4fe;
	16'h2b15 : data <= 32'h832784fe;
	16'h2b16 : data <= 32'h93f7e7ff;
	16'h2b17 : data <= 32'h2324f4fe;
	16'h2b18 : data <= 32'h8327c4fd;
	16'h2b19 : data <= 32'h83a70700;
	16'h2b1a : data <= 32'h032784fe;
	16'h2b1b : data <= 32'h13672700;
	16'h2b1c : data <= 32'h23a2e700;
	16'h2b1d : data <= 32'h6f000003;
	16'h2b1e : data <= 32'h8327c4fd;
	16'h2b1f : data <= 32'h83a70700;
	16'h2b20 : data <= 32'h032784fd;
	16'h2b21 : data <= 32'h03470700;
	16'h2b22 : data <= 32'h23a0e700;
	16'h2b23 : data <= 32'h832784fd;
	16'h2b24 : data <= 32'h93871700;
	16'h2b25 : data <= 32'h232cf4fc;
	16'h2b26 : data <= 32'h832744fd;
	16'h2b27 : data <= 32'h9387f7ff;
	16'h2b28 : data <= 32'h232af4fc;
	16'h2b29 : data <= 32'h832744fd;
	16'h2b2a : data <= 32'h638e0700;
	16'h2b2b : data <= 32'h8327c4fd;
	16'h2b2c : data <= 32'h83a70700;
	16'h2b2d : data <= 32'h83a70701;
	16'h2b2e : data <= 32'h93d7b700;
	16'h2b2f : data <= 32'h93f71700;
	16'h2b30 : data <= 32'he38c07fa;
	16'h2b31 : data <= 32'h8327c4fd;
	16'h2b32 : data <= 32'h032784fd;
	16'h2b33 : data <= 32'h23a2e700;
	16'h2b34 : data <= 32'h8327c4fd;
	16'h2b35 : data <= 32'h032744fd;
	16'h2b36 : data <= 32'h23a4e700;
	16'h2b37 : data <= 32'h8327c4fd;
	16'h2b38 : data <= 32'h032704fd;
	16'h2b39 : data <= 32'h23a6e700;
	16'h2b3a : data <= 32'h6f008002;
	16'h2b3b : data <= 32'h8327c4fd;
	16'h2b3c : data <= 32'h03a70700;
	16'h2b3d : data <= 32'h8327c4fe;
	16'h2b3e : data <= 32'h93861700;
	16'h2b3f : data <= 32'h2326d4fe;
	16'h2b40 : data <= 32'h832684fd;
	16'h2b41 : data <= 32'hb387f600;
	16'h2b42 : data <= 32'h83c70700;
	16'h2b43 : data <= 32'h2320f700;
	16'h2b44 : data <= 32'h0327c4fe;
	16'h2b45 : data <= 32'h832744fd;
	16'h2b46 : data <= 32'h637ef700;
	16'h2b47 : data <= 32'h8327c4fd;
	16'h2b48 : data <= 32'h83a70700;
	16'h2b49 : data <= 32'h83a70701;
	16'h2b4a : data <= 32'h93d7b700;
	16'h2b4b : data <= 32'h93f71700;
	16'h2b4c : data <= 32'he38e07fa;
	16'h2b4d : data <= 32'h8327c4fd;
	16'h2b4e : data <= 32'h13071000;
	16'h2b4f : data <= 32'h23a8e700;
	16'h2b50 : data <= 32'h93070000;
	16'h2b51 : data <= 32'h13850700;
	16'h2b52 : data <= 32'h0324c102;
	16'h2b53 : data <= 32'h13010103;
	16'h2b54 : data <= 32'h67800000;
	16'h2b55 : data <= 32'h130101fd;
	16'h2b56 : data <= 32'h23268102;
	16'h2b57 : data <= 32'h13040103;
	16'h2b58 : data <= 32'h232ea4fc;
	16'h2b59 : data <= 32'h232cb4fc;
	16'h2b5a : data <= 32'h232ac4fc;
	16'h2b5b : data <= 32'h2328d4fc;
	16'h2b5c : data <= 32'h232604fe;
	16'h2b5d : data <= 32'h8327c4fd;
	16'h2b5e : data <= 32'h83a70700;
	16'h2b5f : data <= 32'h83a74700;
	16'h2b60 : data <= 32'h2324f4fe;
	16'h2b61 : data <= 32'h832784fe;
	16'h2b62 : data <= 32'h93f7e7ff;
	16'h2b63 : data <= 32'h2324f4fe;
	16'h2b64 : data <= 32'h8327c4fd;
	16'h2b65 : data <= 32'h83a70700;
	16'h2b66 : data <= 32'h032784fe;
	16'h2b67 : data <= 32'h13672700;
	16'h2b68 : data <= 32'h23a2e700;
	16'h2b69 : data <= 32'h6f004001;
	16'h2b6a : data <= 32'h8327c4fd;
	16'h2b6b : data <= 32'h83a70700;
	16'h2b6c : data <= 32'h83a7c700;
	16'h2b6d : data <= 32'h2322f4fe;
	16'h2b6e : data <= 32'h8327c4fd;
	16'h2b6f : data <= 32'h83a70700;
	16'h2b70 : data <= 32'h83a70701;
	16'h2b71 : data <= 32'h93d77700;
	16'h2b72 : data <= 32'h93f71700;
	16'h2b73 : data <= 32'he38e07fc;
	16'h2b74 : data <= 32'h8327c4fd;
	16'h2b75 : data <= 32'h032784fd;
	16'h2b76 : data <= 32'h23a2e700;
	16'h2b77 : data <= 32'h8327c4fd;
	16'h2b78 : data <= 32'h032744fd;
	16'h2b79 : data <= 32'h23a4e700;
	16'h2b7a : data <= 32'h8327c4fd;
	16'h2b7b : data <= 32'h032704fd;
	16'h2b7c : data <= 32'h23a6e700;
	16'h2b7d : data <= 32'h8327c4fd;
	16'h2b7e : data <= 32'h13072000;
	16'h2b7f : data <= 32'h23a8e700;
	16'h2b80 : data <= 32'h93070000;
	16'h2b81 : data <= 32'h13850700;
	16'h2b82 : data <= 32'h0324c102;
	16'h2b83 : data <= 32'h13010103;
	16'h2b84 : data <= 32'h67800000;
	16'h2b85 : data <= 32'h130101fd;
	16'h2b86 : data <= 32'h23261102;
	16'h2b87 : data <= 32'h23248102;
	16'h2b88 : data <= 32'h13040103;
	16'h2b89 : data <= 32'h232ea4fc;
	16'h2b8a : data <= 32'h8327c4fd;
	16'h2b8b : data <= 32'h03a70701;
	16'h2b8c : data <= 32'h93071000;
	16'h2b8d : data <= 32'h630af700;
	16'h2b8e : data <= 32'h8327c4fd;
	16'h2b8f : data <= 32'h03a70701;
	16'h2b90 : data <= 32'h93072000;
	16'h2b91 : data <= 32'h631cf718;
	16'h2b92 : data <= 32'h8327c4fd;
	16'h2b93 : data <= 32'h83a70700;
	16'h2b94 : data <= 32'h83a70701;
	16'h2b95 : data <= 32'h2326f4fe;
	16'h2b96 : data <= 32'h8327c4fe;
	16'h2b97 : data <= 32'h93f71700;
	16'h2b98 : data <= 32'h63820702;
	16'h2b99 : data <= 32'h8327c4fd;
	16'h2b9a : data <= 32'h13073000;
	16'h2b9b : data <= 32'h23a8e700;
	16'h2b9c : data <= 32'h8327c4fd;
	16'h2b9d : data <= 32'h83a7c700;
	16'h2b9e : data <= 32'h13051003;
	16'h2b9f : data <= 32'he7800700;
	16'h2ba0 : data <= 32'h6f000016;
	16'h2ba1 : data <= 32'h8327c4fe;
	16'h2ba2 : data <= 32'h93d73700;
	16'h2ba3 : data <= 32'h93f71700;
	16'h2ba4 : data <= 32'h63820702;
	16'h2ba5 : data <= 32'h8327c4fd;
	16'h2ba6 : data <= 32'h13073000;
	16'h2ba7 : data <= 32'h23a8e700;
	16'h2ba8 : data <= 32'h8327c4fd;
	16'h2ba9 : data <= 32'h83a7c700;
	16'h2baa : data <= 32'h13052003;
	16'h2bab : data <= 32'he7800700;
	16'h2bac : data <= 32'h6f000013;
	16'h2bad : data <= 32'h8327c4fe;
	16'h2bae : data <= 32'h93d72700;
	16'h2baf : data <= 32'h93f71700;
	16'h2bb0 : data <= 32'h63820702;
	16'h2bb1 : data <= 32'h8327c4fd;
	16'h2bb2 : data <= 32'h13073000;
	16'h2bb3 : data <= 32'h23a8e700;
	16'h2bb4 : data <= 32'h8327c4fd;
	16'h2bb5 : data <= 32'h83a7c700;
	16'h2bb6 : data <= 32'h13050000;
	16'h2bb7 : data <= 32'he7800700;
	16'h2bb8 : data <= 32'h6f000010;
	16'h2bb9 : data <= 32'h8327c4fd;
	16'h2bba : data <= 32'h03a70701;
	16'h2bbb : data <= 32'h93071000;
	16'h2bbc : data <= 32'h6316f70c;
	16'h2bbd : data <= 32'h6f004005;
	16'h2bbe : data <= 32'h8327c4fd;
	16'h2bbf : data <= 32'h83a70700;
	16'h2bc0 : data <= 32'h0327c4fd;
	16'h2bc1 : data <= 32'h03274700;
	16'h2bc2 : data <= 32'h03470700;
	16'h2bc3 : data <= 32'h23a0e700;
	16'h2bc4 : data <= 32'h8327c4fd;
	16'h2bc5 : data <= 32'h83a74700;
	16'h2bc6 : data <= 32'h13871700;
	16'h2bc7 : data <= 32'h8327c4fd;
	16'h2bc8 : data <= 32'h23a2e700;
	16'h2bc9 : data <= 32'h8327c4fd;
	16'h2bca : data <= 32'h83a78700;
	16'h2bcb : data <= 32'h1387f7ff;
	16'h2bcc : data <= 32'h8327c4fd;
	16'h2bcd : data <= 32'h23a4e700;
	16'h2bce : data <= 32'h8327c4fd;
	16'h2bcf : data <= 32'h83a70700;
	16'h2bd0 : data <= 32'h83a70701;
	16'h2bd1 : data <= 32'h2326f4fe;
	16'h2bd2 : data <= 32'h8327c4fe;
	16'h2bd3 : data <= 32'h93d7b700;
	16'h2bd4 : data <= 32'h93f71700;
	16'h2bd5 : data <= 32'h63960708;
	16'h2bd6 : data <= 32'h8327c4fd;
	16'h2bd7 : data <= 32'h83a78700;
	16'h2bd8 : data <= 32'he39c07f8;
	16'h2bd9 : data <= 32'h6f00c007;
	16'h2bda : data <= 32'h8327c4fd;
	16'h2bdb : data <= 32'h83a74700;
	16'h2bdc : data <= 32'h0327c4fd;
	16'h2bdd : data <= 32'h03270700;
	16'h2bde : data <= 32'h0327c700;
	16'h2bdf : data <= 32'h1377f70f;
	16'h2be0 : data <= 32'h2380e700;
	16'h2be1 : data <= 32'h8327c4fd;
	16'h2be2 : data <= 32'h83a74700;
	16'h2be3 : data <= 32'h13871700;
	16'h2be4 : data <= 32'h8327c4fd;
	16'h2be5 : data <= 32'h23a2e700;
	16'h2be6 : data <= 32'h8327c4fd;
	16'h2be7 : data <= 32'h83a78700;
	16'h2be8 : data <= 32'h1387f7ff;
	16'h2be9 : data <= 32'h8327c4fd;
	16'h2bea : data <= 32'h23a4e700;
	16'h2beb : data <= 32'h8327c4fd;
	16'h2bec : data <= 32'h83a70700;
	16'h2bed : data <= 32'h83a70701;
	16'h2bee : data <= 32'h2326f4fe;
	16'h2bef : data <= 32'h8327c4fe;
	16'h2bf0 : data <= 32'h93d77700;
	16'h2bf1 : data <= 32'h93f71700;
	16'h2bf2 : data <= 32'h639c0700;
	16'h2bf3 : data <= 32'h8327c4fd;
	16'h2bf4 : data <= 32'h83a78700;
	16'h2bf5 : data <= 32'he39a07f8;
	16'h2bf6 : data <= 32'h6f008000;
	16'h2bf7 : data <= 32'h13000000;
	16'h2bf8 : data <= 32'h8320c102;
	16'h2bf9 : data <= 32'h03248102;
	16'h2bfa : data <= 32'h13010103;
	16'h2bfb : data <= 32'h67800000;
	16'h2bfc : data <= 32'h130101fc;
	16'h2bfd : data <= 32'h232e8102;
	16'h2bfe : data <= 32'h13040104;
	16'h2bff : data <= 32'h2326a4fc;
	16'h2c00 : data <= 32'h2324b4fc;
	16'h2c01 : data <= 32'h2322c4fc;
	16'h2c02 : data <= 32'h2320d4fc;
	16'h2c03 : data <= 32'h232604fe;
	16'h2c04 : data <= 32'h032744fc;
	16'h2c05 : data <= 32'h93070004;
	16'h2c06 : data <= 32'h63f6e700;
	16'h2c07 : data <= 32'h93070003;
	16'h2c08 : data <= 32'h6f004016;
	16'h2c09 : data <= 32'h032744fc;
	16'h2c0a : data <= 32'h93070004;
	16'h2c0b : data <= 32'h631af702;
	16'h2c0c : data <= 32'h8327c4fc;
	16'h2c0d : data <= 32'h83a70700;
	16'h2c0e : data <= 32'h83a74700;
	16'h2c0f : data <= 32'h2324f4fe;
	16'h2c10 : data <= 32'h832784fe;
	16'h2c11 : data <= 32'h93f707fc;
	16'h2c12 : data <= 32'h2324f4fe;
	16'h2c13 : data <= 32'h8327c4fc;
	16'h2c14 : data <= 32'h83a70700;
	16'h2c15 : data <= 32'h032784fe;
	16'h2c16 : data <= 32'h23a2e700;
	16'h2c17 : data <= 32'h6f000004;
	16'h2c18 : data <= 32'h8327c4fc;
	16'h2c19 : data <= 32'h83a70700;
	16'h2c1a : data <= 32'h83a74700;
	16'h2c1b : data <= 32'h2322f4fe;
	16'h2c1c : data <= 32'h832744fe;
	16'h2c1d : data <= 32'h93f707fc;
	16'h2c1e : data <= 32'h2322f4fe;
	16'h2c1f : data <= 32'h8327c4fc;
	16'h2c20 : data <= 32'h83a70700;
	16'h2c21 : data <= 32'h032744fc;
	16'h2c22 : data <= 32'h13172700;
	16'h2c23 : data <= 32'h9376f70f;
	16'h2c24 : data <= 32'h032744fe;
	16'h2c25 : data <= 32'h33e7e600;
	16'h2c26 : data <= 32'h23a2e700;
	16'h2c27 : data <= 32'h8327c4fc;
	16'h2c28 : data <= 32'h83a70700;
	16'h2c29 : data <= 32'h83a74700;
	16'h2c2a : data <= 32'h2320f4fe;
	16'h2c2b : data <= 32'h832704fe;
	16'h2c2c : data <= 32'h93f7e7ff;
	16'h2c2d : data <= 32'h2320f4fe;
	16'h2c2e : data <= 32'h8327c4fc;
	16'h2c2f : data <= 32'h83a70700;
	16'h2c30 : data <= 32'h032704fe;
	16'h2c31 : data <= 32'h23a2e700;
	16'h2c32 : data <= 32'h8327c4fc;
	16'h2c33 : data <= 32'h83a70700;
	16'h2c34 : data <= 32'h83a74700;
	16'h2c35 : data <= 32'h232ef4fc;
	16'h2c36 : data <= 32'h8327c4fd;
	16'h2c37 : data <= 32'h93f7e7ff;
	16'h2c38 : data <= 32'h232ef4fc;
	16'h2c39 : data <= 32'h8327c4fc;
	16'h2c3a : data <= 32'h83a70700;
	16'h2c3b : data <= 32'h0327c4fd;
	16'h2c3c : data <= 32'h23a2e700;
	16'h2c3d : data <= 32'h6f004001;
	16'h2c3e : data <= 32'h8327c4fc;
	16'h2c3f : data <= 32'h83a70700;
	16'h2c40 : data <= 32'h83a7c700;
	16'h2c41 : data <= 32'h232cf4fc;
	16'h2c42 : data <= 32'h8327c4fc;
	16'h2c43 : data <= 32'h83a70700;
	16'h2c44 : data <= 32'h83a70701;
	16'h2c45 : data <= 32'h93d77700;
	16'h2c46 : data <= 32'h93f71700;
	16'h2c47 : data <= 32'he38e07fc;
	16'h2c48 : data <= 32'h8327c4fc;
	16'h2c49 : data <= 32'h032784fc;
	16'h2c4a : data <= 32'h23a2e700;
	16'h2c4b : data <= 32'h8327c4fc;
	16'h2c4c : data <= 32'h032744fc;
	16'h2c4d : data <= 32'h23a4e700;
	16'h2c4e : data <= 32'h8327c4fc;
	16'h2c4f : data <= 32'h032704fc;
	16'h2c50 : data <= 32'h23a6e700;
	16'h2c51 : data <= 32'h8327c4fc;
	16'h2c52 : data <= 32'h83a70700;
	16'h2c53 : data <= 32'h83a74700;
	16'h2c54 : data <= 32'h232af4fc;
	16'h2c55 : data <= 32'h832744fd;
	16'h2c56 : data <= 32'h93f7e7ff;
	16'h2c57 : data <= 32'h232af4fc;
	16'h2c58 : data <= 32'h8327c4fc;
	16'h2c59 : data <= 32'h83a70700;
	16'h2c5a : data <= 32'h032744fd;
	16'h2c5b : data <= 32'h13670720;
	16'h2c5c : data <= 32'h23a2e700;
	16'h2c5d : data <= 32'h8327c4fc;
	16'h2c5e : data <= 32'h13072000;
	16'h2c5f : data <= 32'h23a8e700;
	16'h2c60 : data <= 32'h93070000;
	16'h2c61 : data <= 32'h13850700;
	16'h2c62 : data <= 32'h0324c103;
	16'h2c63 : data <= 32'h13010104;
	16'h2c64 : data <= 32'h67800000;
	16'h2c65 : data <= 32'h130101fd;
	16'h2c66 : data <= 32'h23268102;
	16'h2c67 : data <= 32'h13040103;
	16'h2c68 : data <= 32'h232ea4fc;
	16'h2c69 : data <= 32'h232cb4fc;
	16'h2c6a : data <= 32'h232ac4fc;
	16'h2c6b : data <= 32'h232604fe;
	16'h2c6c : data <= 32'h232604fe;
	16'h2c6d : data <= 32'h6f008004;
	16'h2c6e : data <= 32'h13000000;
	16'h2c6f : data <= 32'h8327c4fd;
	16'h2c70 : data <= 32'h83a70700;
	16'h2c71 : data <= 32'h83a7c700;
	16'h2c72 : data <= 32'h93d72700;
	16'h2c73 : data <= 32'h93f71700;
	16'h2c74 : data <= 32'he39607fe;
	16'h2c75 : data <= 32'h8327c4fd;
	16'h2c76 : data <= 32'h83a70700;
	16'h2c77 : data <= 32'h0327c4fe;
	16'h2c78 : data <= 32'h832684fd;
	16'h2c79 : data <= 32'h3387e600;
	16'h2c7a : data <= 32'h03470700;
	16'h2c7b : data <= 32'h23a2e700;
	16'h2c7c : data <= 32'h8327c4fe;
	16'h2c7d : data <= 32'h93871700;
	16'h2c7e : data <= 32'h2326f4fe;
	16'h2c7f : data <= 32'h0327c4fe;
	16'h2c80 : data <= 32'h832744fd;
	16'h2c81 : data <= 32'he36af7fa;
	16'h2c82 : data <= 32'h93070000;
	16'h2c83 : data <= 32'h13850700;
	16'h2c84 : data <= 32'h0324c102;
	16'h2c85 : data <= 32'h13010103;
	16'h2c86 : data <= 32'h67800000;
	16'h2c87 : data <= 32'h130101fd;
	16'h2c88 : data <= 32'h23268102;
	16'h2c89 : data <= 32'h13040103;
	16'h2c8a : data <= 32'h232ea4fc;
	16'h2c8b : data <= 32'h232cb4fc;
	16'h2c8c : data <= 32'h232ac4fc;
	16'h2c8d : data <= 32'h232604fe;
	16'h2c8e : data <= 32'h232604fe;
	16'h2c8f : data <= 32'h6f00c004;
	16'h2c90 : data <= 32'h13000000;
	16'h2c91 : data <= 32'h8327c4fd;
	16'h2c92 : data <= 32'h83a70700;
	16'h2c93 : data <= 32'h83a7c700;
	16'h2c94 : data <= 32'h93d75700;
	16'h2c95 : data <= 32'h93f71700;
	16'h2c96 : data <= 32'he39607fe;
	16'h2c97 : data <= 32'h8327c4fe;
	16'h2c98 : data <= 32'h032784fd;
	16'h2c99 : data <= 32'hb307f700;
	16'h2c9a : data <= 32'h0327c4fd;
	16'h2c9b : data <= 32'h03270700;
	16'h2c9c : data <= 32'h03278700;
	16'h2c9d : data <= 32'h1377f70f;
	16'h2c9e : data <= 32'h2380e700;
	16'h2c9f : data <= 32'h8327c4fe;
	16'h2ca0 : data <= 32'h93871700;
	16'h2ca1 : data <= 32'h2326f4fe;
	16'h2ca2 : data <= 32'h0327c4fe;
	16'h2ca3 : data <= 32'h832744fd;
	16'h2ca4 : data <= 32'he368f7fa;
	16'h2ca5 : data <= 32'h93070000;
	16'h2ca6 : data <= 32'h13850700;
	16'h2ca7 : data <= 32'h0324c102;
	16'h2ca8 : data <= 32'h13010103;
	16'h2ca9 : data <= 32'h67800000;
	16'h2caa : data <= 32'h130101fe;
	16'h2cab : data <= 32'h232e1100;
	16'h2cac : data <= 32'h232c8100;
	16'h2cad : data <= 32'h13040102;
	16'h2cae : data <= 32'h2326a4fe;
	16'h2caf : data <= 32'h2324b4fe;
	16'h2cb0 : data <= 32'h2322c4fe;
	16'h2cb1 : data <= 32'h2320d4fe;
	16'h2cb2 : data <= 32'h8327c4fe;
	16'h2cb3 : data <= 32'h83a70702;
	16'h2cb4 : data <= 32'h63960700;
	16'h2cb5 : data <= 32'h93070002;
	16'h2cb6 : data <= 32'h6f00c00c;
	16'h2cb7 : data <= 32'h8327c4fe;
	16'h2cb8 : data <= 32'h03a70702;
	16'h2cb9 : data <= 32'h93071000;
	16'h2cba : data <= 32'h6316f700;
	16'h2cbb : data <= 32'h93071002;
	16'h2cbc : data <= 32'h6f00400b;
	16'h2cbd : data <= 32'h8327c4fe;
	16'h2cbe : data <= 32'h03a70702;
	16'h2cbf : data <= 32'h93072000;
	16'h2cc0 : data <= 32'h630cf702;
	16'h2cc1 : data <= 32'h93071000;
	16'h2cc2 : data <= 32'h6f00c009;
	16'h2cc3 : data <= 32'h8327c4fe;
	16'h2cc4 : data <= 32'h83a70700;
	16'h2cc5 : data <= 32'h032784fe;
	16'h2cc6 : data <= 32'h03470700;
	16'h2cc7 : data <= 32'h23a2e700;
	16'h2cc8 : data <= 32'h832784fe;
	16'h2cc9 : data <= 32'h93871700;
	16'h2cca : data <= 32'h2324f4fe;
	16'h2ccb : data <= 32'h832744fe;
	16'h2ccc : data <= 32'h9387f7ff;
	16'h2ccd : data <= 32'h2322f4fe;
	16'h2cce : data <= 32'h832744fe;
	16'h2ccf : data <= 32'h638e0700;
	16'h2cd0 : data <= 32'h8327c4fe;
	16'h2cd1 : data <= 32'h83a70700;
	16'h2cd2 : data <= 32'h83a7c700;
	16'h2cd3 : data <= 32'h93d72700;
	16'h2cd4 : data <= 32'h93f71700;
	16'h2cd5 : data <= 32'he38c07fa;
	16'h2cd6 : data <= 32'h832744fe;
	16'h2cd7 : data <= 32'h639a0700;
	16'h2cd8 : data <= 32'h832704fe;
	16'h2cd9 : data <= 32'he7800700;
	16'h2cda : data <= 32'h93070000;
	16'h2cdb : data <= 32'h6f008003;
	16'h2cdc : data <= 32'h8327c4fe;
	16'h2cdd : data <= 32'h032784fe;
	16'h2cde : data <= 32'h23a2e700;
	16'h2cdf : data <= 32'h8327c4fe;
	16'h2ce0 : data <= 32'h032744fe;
	16'h2ce1 : data <= 32'h23a6e700;
	16'h2ce2 : data <= 32'h8327c4fe;
	16'h2ce3 : data <= 32'h032704fe;
	16'h2ce4 : data <= 32'h23aae700;
	16'h2ce5 : data <= 32'h8327c4fe;
	16'h2ce6 : data <= 32'h13071000;
	16'h2ce7 : data <= 32'h23a0e702;
	16'h2ce8 : data <= 32'h93070000;
	16'h2ce9 : data <= 32'h13850700;
	16'h2cea : data <= 32'h8320c101;
	16'h2ceb : data <= 32'h03248101;
	16'h2cec : data <= 32'h13010102;
	16'h2ced : data <= 32'h67800000;
	16'h2cee : data <= 32'h130101fe;
	16'h2cef : data <= 32'h232e1100;
	16'h2cf0 : data <= 32'h232c8100;
	16'h2cf1 : data <= 32'h13040102;
	16'h2cf2 : data <= 32'h2326a4fe;
	16'h2cf3 : data <= 32'h2324b4fe;
	16'h2cf4 : data <= 32'h93070600;
	16'h2cf5 : data <= 32'h2320d4fe;
	16'h2cf6 : data <= 32'h2313f4fe;
	16'h2cf7 : data <= 32'h8327c4fe;
	16'h2cf8 : data <= 32'h83a70702;
	16'h2cf9 : data <= 32'h63960700;
	16'h2cfa : data <= 32'h93070002;
	16'h2cfb : data <= 32'h6f00000d;
	16'h2cfc : data <= 32'h8327c4fe;
	16'h2cfd : data <= 32'h03a70702;
	16'h2cfe : data <= 32'h93071000;
	16'h2cff : data <= 32'h6316f700;
	16'h2d00 : data <= 32'h93071002;
	16'h2d01 : data <= 32'h6f00800b;
	16'h2d02 : data <= 32'h8327c4fe;
	16'h2d03 : data <= 32'h03a70702;
	16'h2d04 : data <= 32'h93072000;
	16'h2d05 : data <= 32'h630ef702;
	16'h2d06 : data <= 32'h93071000;
	16'h2d07 : data <= 32'h6f00000a;
	16'h2d08 : data <= 32'h8327c4fe;
	16'h2d09 : data <= 32'h83a70700;
	16'h2d0a : data <= 32'h83a78700;
	16'h2d0b : data <= 32'h13f7f70f;
	16'h2d0c : data <= 32'h832784fe;
	16'h2d0d : data <= 32'h2380e700;
	16'h2d0e : data <= 32'h832784fe;
	16'h2d0f : data <= 32'h93871700;
	16'h2d10 : data <= 32'h2324f4fe;
	16'h2d11 : data <= 32'h835764fe;
	16'h2d12 : data <= 32'h9387f7ff;
	16'h2d13 : data <= 32'h2313f4fe;
	16'h2d14 : data <= 32'h835764fe;
	16'h2d15 : data <= 32'h638e0700;
	16'h2d16 : data <= 32'h8327c4fe;
	16'h2d17 : data <= 32'h83a70700;
	16'h2d18 : data <= 32'h83a7c700;
	16'h2d19 : data <= 32'h93d75700;
	16'h2d1a : data <= 32'h93f71700;
	16'h2d1b : data <= 32'he38a07fa;
	16'h2d1c : data <= 32'h835764fe;
	16'h2d1d : data <= 32'h639a0700;
	16'h2d1e : data <= 32'h832704fe;
	16'h2d1f : data <= 32'he7800700;
	16'h2d20 : data <= 32'h93070000;
	16'h2d21 : data <= 32'h6f008003;
	16'h2d22 : data <= 32'h8327c4fe;
	16'h2d23 : data <= 32'h032784fe;
	16'h2d24 : data <= 32'h23a4e700;
	16'h2d25 : data <= 32'h035764fe;
	16'h2d26 : data <= 32'h8327c4fe;
	16'h2d27 : data <= 32'h23a8e700;
	16'h2d28 : data <= 32'h8327c4fe;
	16'h2d29 : data <= 32'h032704fe;
	16'h2d2a : data <= 32'h23ace700;
	16'h2d2b : data <= 32'h8327c4fe;
	16'h2d2c : data <= 32'h13071000;
	16'h2d2d : data <= 32'h23aee700;
	16'h2d2e : data <= 32'h93070000;
	16'h2d2f : data <= 32'h13850700;
	16'h2d30 : data <= 32'h8320c101;
	16'h2d31 : data <= 32'h03248101;
	16'h2d32 : data <= 32'h13010102;
	16'h2d33 : data <= 32'h67800000;
	16'h2d34 : data <= 32'h130101fd;
	16'h2d35 : data <= 32'h23261102;
	16'h2d36 : data <= 32'h23248102;
	16'h2d37 : data <= 32'h13040103;
	16'h2d38 : data <= 32'h232ea4fc;
	16'h2d39 : data <= 32'h8327c4fd;
	16'h2d3a : data <= 32'h03a70702;
	16'h2d3b : data <= 32'h93071000;
	16'h2d3c : data <= 32'h6316f70a;
	16'h2d3d : data <= 32'h8327c4fd;
	16'h2d3e : data <= 32'h83a7c700;
	16'h2d3f : data <= 32'h2326f4fe;
	16'h2d40 : data <= 32'h6f004004;
	16'h2d41 : data <= 32'h8327c4fd;
	16'h2d42 : data <= 32'h83a70700;
	16'h2d43 : data <= 32'h0327c4fd;
	16'h2d44 : data <= 32'h03274700;
	16'h2d45 : data <= 32'h03470700;
	16'h2d46 : data <= 32'h23a2e700;
	16'h2d47 : data <= 32'h8327c4fd;
	16'h2d48 : data <= 32'h83a74700;
	16'h2d49 : data <= 32'h13871700;
	16'h2d4a : data <= 32'h8327c4fd;
	16'h2d4b : data <= 32'h23a2e700;
	16'h2d4c : data <= 32'h8327c4fd;
	16'h2d4d : data <= 32'h83a7c700;
	16'h2d4e : data <= 32'h1387f7ff;
	16'h2d4f : data <= 32'h8327c4fd;
	16'h2d50 : data <= 32'h23a6e700;
	16'h2d51 : data <= 32'h8327c4fd;
	16'h2d52 : data <= 32'h83a7c700;
	16'h2d53 : data <= 32'h638e0700;
	16'h2d54 : data <= 32'h8327c4fd;
	16'h2d55 : data <= 32'h83a70700;
	16'h2d56 : data <= 32'h83a7c700;
	16'h2d57 : data <= 32'h93d72700;
	16'h2d58 : data <= 32'h93f71700;
	16'h2d59 : data <= 32'he38007fa;
	16'h2d5a : data <= 32'h8327c4fd;
	16'h2d5b : data <= 32'h83a7c700;
	16'h2d5c : data <= 32'h639a0702;
	16'h2d5d : data <= 32'h8327c4fe;
	16'h2d5e : data <= 32'h63860702;
	16'h2d5f : data <= 32'h8327c4fd;
	16'h2d60 : data <= 32'h83a74701;
	16'h2d61 : data <= 32'he7800700;
	16'h2d62 : data <= 32'h8327c4fd;
	16'h2d63 : data <= 32'h13072000;
	16'h2d64 : data <= 32'h23a0e702;
	16'h2d65 : data <= 32'h13000000;
	16'h2d66 : data <= 32'h6f00c000;
	16'h2d67 : data <= 32'h13000000;
	16'h2d68 : data <= 32'h6f008000;
	16'h2d69 : data <= 32'h13000000;
	16'h2d6a : data <= 32'h8320c102;
	16'h2d6b : data <= 32'h03248102;
	16'h2d6c : data <= 32'h13010103;
	16'h2d6d : data <= 32'h67800000;
	16'h2d6e : data <= 32'h130101fd;
	16'h2d6f : data <= 32'h23261102;
	16'h2d70 : data <= 32'h23248102;
	16'h2d71 : data <= 32'h13040103;
	16'h2d72 : data <= 32'h232ea4fc;
	16'h2d73 : data <= 32'h8327c4fd;
	16'h2d74 : data <= 32'h03a7c701;
	16'h2d75 : data <= 32'h93071000;
	16'h2d76 : data <= 32'h6318f70a;
	16'h2d77 : data <= 32'h8327c4fd;
	16'h2d78 : data <= 32'h83a70701;
	16'h2d79 : data <= 32'h2326f4fe;
	16'h2d7a : data <= 32'h6f008004;
	16'h2d7b : data <= 32'h8327c4fd;
	16'h2d7c : data <= 32'h83a78700;
	16'h2d7d : data <= 32'h0327c4fd;
	16'h2d7e : data <= 32'h03270700;
	16'h2d7f : data <= 32'h03278700;
	16'h2d80 : data <= 32'h1377f70f;
	16'h2d81 : data <= 32'h2380e700;
	16'h2d82 : data <= 32'h8327c4fd;
	16'h2d83 : data <= 32'h83a78700;
	16'h2d84 : data <= 32'h13871700;
	16'h2d85 : data <= 32'h8327c4fd;
	16'h2d86 : data <= 32'h23a4e700;
	16'h2d87 : data <= 32'h8327c4fd;
	16'h2d88 : data <= 32'h83a70701;
	16'h2d89 : data <= 32'h1387f7ff;
	16'h2d8a : data <= 32'h8327c4fd;
	16'h2d8b : data <= 32'h23a8e700;
	16'h2d8c : data <= 32'h8327c4fd;
	16'h2d8d : data <= 32'h83a70701;
	16'h2d8e : data <= 32'h638e0700;
	16'h2d8f : data <= 32'h8327c4fd;
	16'h2d90 : data <= 32'h83a70700;
	16'h2d91 : data <= 32'h83a7c700;
	16'h2d92 : data <= 32'h93d75700;
	16'h2d93 : data <= 32'h93f71700;
	16'h2d94 : data <= 32'he38e07f8;
	16'h2d95 : data <= 32'h8327c4fd;
	16'h2d96 : data <= 32'h83a70701;
	16'h2d97 : data <= 32'h639a0702;
	16'h2d98 : data <= 32'h8327c4fe;
	16'h2d99 : data <= 32'h63860702;
	16'h2d9a : data <= 32'h8327c4fd;
	16'h2d9b : data <= 32'h83a78701;
	16'h2d9c : data <= 32'he7800700;
	16'h2d9d : data <= 32'h8327c4fd;
	16'h2d9e : data <= 32'h13072000;
	16'h2d9f : data <= 32'h23aee700;
	16'h2da0 : data <= 32'h13000000;
	16'h2da1 : data <= 32'h6f00c000;
	16'h2da2 : data <= 32'h13000000;
	16'h2da3 : data <= 32'h6f008000;
	16'h2da4 : data <= 32'h13000000;
	16'h2da5 : data <= 32'h8320c102;
	16'h2da6 : data <= 32'h03248102;
	16'h2da7 : data <= 32'h13010103;
	16'h2da8 : data <= 32'h67800000;
	16'h2da9 : data <= 32'h4743433a;
	16'h2daa : data <= 32'h2028474e;
	16'h2dab : data <= 32'h55292035;
	16'h2dac : data <= 32'h2e332e30;
	16'h2dad : data <= 32'h00800080;
	16'h2dae : data <= 32'h02000000;
	16'h2daf : data <= 32'h02000000;
	16'h2db0 : data <= 32'h00100080;
	16'h2db1 : data <= 32'h03000000;
	16'h2db2 : data <= 32'hFF;
	default : data <= 32'hDEADBEEF;
	//default : data <= 32'b0;
endcase 
end 
else begin data <= TOPRAMdata; end
 end
 always_comb begin  if(addr >= 16'h2db3) begin topw_en = w_en; end else begin topw_en = 0; end end endmodule
