VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO dig_poly_NAND_NOR2_x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN dig_poly_NAND_NOR2_x1 0 0 ;
  SIZE 10.25 BY 2.56 ;
  SYMMETRY X Y ;
  SITE CoreSite8T ;
  PIN orient
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.915 0.66 1.135 1.58 ;
      LAYER M1 ;
        RECT 0.935 0.99 1.115 1.21 ;
        RECT 0.945 0.66 1.105 1.58 ;
      LAYER V12 ;
        RECT 0.955 1.03 1.095 1.17 ;
    END
  END orient
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.335 1.57 6.105 1.73 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.605 1.535 7.155 1.775 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.675 1.96 7.485 2.16 ;
        RECT 7.325 0.47 7.485 2.16 ;
        RECT 6.675 1.16 7.485 1.36 ;
        RECT 6.675 0.47 7.485 0.67 ;
    END
  END X
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.33 10.25 2.56 ;
        RECT 3.815 1.54 3.975 2.56 ;
        RECT 2.995 2.06 3.155 2.56 ;
        RECT 2.175 1.54 2.335 2.56 ;
        RECT 1.765 1.54 1.925 2.56 ;
        RECT 0.945 2.06 1.105 2.56 ;
        RECT 0.125 1.54 0.285 2.56 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 10.25 0.23 ;
        RECT 3.815 0 3.975 0.76 ;
        RECT 2.995 0 3.155 0.5 ;
        RECT 2.175 0 2.335 0.76 ;
        RECT 1.765 0 1.925 0.76 ;
        RECT 0.945 0 1.105 0.5 ;
        RECT 0.125 0 0.285 0.76 ;
    END
  END vss!
  OBS
    LAYER M1 ;
      RECT 8.69 1.97 8.955 2.17 ;
      RECT 8.775 0.39 8.955 2.17 ;
      RECT 7.645 1.97 8.44 2.17 ;
      RECT 7.645 1.16 7.805 2.17 ;
      RECT 7.965 1.21 8.205 1.41 ;
      RECT 7.965 0.86 8.105 1.41 ;
      RECT 7.645 0.86 8.105 1 ;
      RECT 7.645 0.47 7.805 1 ;
      RECT 5.865 1.21 6.105 1.41 ;
      RECT 5.965 0.86 6.105 1.41 ;
      RECT 5.965 0.86 6.415 1 ;
      RECT 6.265 0.47 6.415 1 ;
      RECT 6.265 0.47 6.425 0.67 ;
      RECT 5.25 1.96 6.425 2.17 ;
      RECT 6.265 1.16 6.425 2.17 ;
      RECT 4.84 0.755 5 2.17 ;
      RECT 4.84 0.755 5.295 0.975 ;
      RECT 5.115 0.39 5.295 0.975 ;
      RECT 3.395 0.39 3.575 2.13 ;
      RECT 2.585 0.39 2.745 2.13 ;
      RECT 2.585 1.74 3.575 1.9 ;
      RECT 2.575 1.66 2.755 1.88 ;
      RECT 2.995 0.66 3.155 1.58 ;
      RECT 2.985 0.99 3.165 1.21 ;
      RECT 1.345 0.39 1.525 2.14 ;
      RECT 0.535 0.39 0.695 2.13 ;
      RECT 0.535 1.74 1.525 1.9 ;
      RECT 9.115 1.71 9.335 2.17 ;
      RECT 8.455 0.42 8.615 1.41 ;
      RECT 7.965 0.39 8.295 0.7 ;
      RECT 5.775 0.39 6.105 0.7 ;
      RECT 5.455 0.42 5.615 1.41 ;
      RECT 4.46 1.71 4.68 2.17 ;
    LAYER V12 ;
      RECT 9.155 2.01 9.295 2.15 ;
      RECT 8.795 0.795 8.935 0.935 ;
      RECT 8.055 0.52 8.195 0.66 ;
      RECT 5.875 0.52 6.015 0.66 ;
      RECT 5.135 0.795 5.275 0.935 ;
      RECT 4.5 2.01 4.64 2.15 ;
      RECT 3.415 0.46 3.555 0.6 ;
      RECT 3.415 0.74 3.555 0.88 ;
      RECT 3.415 1.42 3.555 1.56 ;
      RECT 3.415 1.7 3.555 1.84 ;
      RECT 3.005 1.03 3.145 1.17 ;
      RECT 2.595 1.7 2.735 1.84 ;
      RECT 1.365 0.46 1.505 0.6 ;
      RECT 1.365 0.74 1.505 0.88 ;
      RECT 1.365 1.4 1.505 1.54 ;
      RECT 1.365 1.68 1.505 1.82 ;
      RECT 1.365 1.96 1.505 2.1 ;
    LAYER M2 ;
      RECT 1.325 2.17 9.315 2.4 ;
      RECT 9.135 1.97 9.315 2.4 ;
      RECT 7.53 0.5 7.71 2.4 ;
      RECT 4.48 1.97 4.66 2.4 ;
      RECT 1.325 0.39 1.545 2.4 ;
      RECT 2.965 0.66 3.185 1.58 ;
      RECT 1.325 0.66 3.185 0.89 ;
      RECT 8.015 0.5 8.235 0.68 ;
      RECT 5.835 0.5 6.055 0.68 ;
      RECT 5.835 0.5 8.235 0.66 ;
      RECT 2.555 1.74 3.595 1.92 ;
      RECT 3.375 0.16 3.595 1.92 ;
      RECT 2.555 1.68 2.775 1.92 ;
      RECT 8.425 0.775 8.975 0.955 ;
      RECT 5.095 0.775 5.645 0.955 ;
      RECT 5.425 0.16 5.645 0.955 ;
      RECT 8.425 0.155 8.645 0.955 ;
      RECT 3.375 0.16 8.645 0.34 ;
  END
END dig_poly_NAND_NOR2_x1

MACRO dig_poly_XOR_BUF2_x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN dig_poly_XOR_BUF2_x1 0 0 ;
  SIZE 14.35 BY 2.56 ;
  SYMMETRY X Y ;
  SITE CoreSite8T ;
  PIN orient
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.945 0.66 1.105 1.58 ;
    END
  END orient
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 13.47 1.735 14.12 2.03 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 13.47 0.53 14.115 0.87 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.085 1.595 12.265 1.815 ;
        RECT 12.105 1.2 12.245 1.815 ;
        RECT 7.59 1.2 12.245 1.34 ;
        RECT 11.675 0.775 11.855 0.995 ;
        RECT 11.695 0.775 11.835 1.34 ;
        RECT 10.235 1.595 10.415 1.815 ;
        RECT 10.255 1.2 10.395 1.815 ;
        RECT 7.59 1.18 7.81 1.36 ;
      LAYER M1 ;
        RECT 12.005 1.54 12.455 1.81 ;
        RECT 11.62 0.515 11.93 0.99 ;
        RECT 10.165 1.555 10.595 1.82 ;
        RECT 7.425 1.605 7.8 1.805 ;
        RECT 7.6 0.785 7.8 1.805 ;
        RECT 7.445 0.785 7.8 0.985 ;
      LAYER V12 ;
        RECT 7.63 1.2 7.77 1.34 ;
        RECT 10.255 1.635 10.395 1.775 ;
        RECT 11.695 0.815 11.835 0.955 ;
        RECT 12.105 1.635 12.245 1.775 ;
    END
  END X
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.33 14.35 2.56 ;
        RECT 3.815 1.54 3.975 2.56 ;
        RECT 2.995 2.06 3.155 2.56 ;
        RECT 2.175 1.54 2.335 2.56 ;
        RECT 1.765 1.54 1.925 2.56 ;
        RECT 0.945 2.06 1.105 2.56 ;
        RECT 0.125 1.54 0.285 2.56 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 14.35 0.23 ;
        RECT 3.815 0 3.975 0.76 ;
        RECT 2.995 0 3.155 0.5 ;
        RECT 2.175 0 2.335 0.76 ;
        RECT 1.765 0 1.925 0.76 ;
        RECT 0.945 0 1.105 0.5 ;
        RECT 0.125 0 0.285 0.76 ;
    END
  END vss!
  OBS
    LAYER M1 ;
      RECT 13.025 0.785 13.185 1.805 ;
      RECT 12.995 0.795 13.215 0.975 ;
      RECT 12.17 1.985 12.88 2.165 ;
      RECT 12.335 1.97 12.555 2.165 ;
      RECT 12.615 1.22 12.775 1.805 ;
      RECT 11.165 1.22 12.775 1.38 ;
      RECT 11.165 0.785 11.325 1.38 ;
      RECT 9.565 1.97 9.785 2.15 ;
      RECT 9.565 1.98 10.915 2.14 ;
      RECT 10.755 0.785 10.915 2.14 ;
      RECT 9.31 1.97 9.785 2.13 ;
      RECT 9.31 1.605 9.47 2.13 ;
      RECT 9.835 1.225 9.995 1.805 ;
      RECT 9.835 1.225 10.405 1.385 ;
      RECT 10.245 0.785 10.405 1.385 ;
      RECT 9.31 0.785 9.995 0.985 ;
      RECT 7.035 0.395 7.195 0.985 ;
      RECT 9.31 0.395 9.47 0.985 ;
      RECT 7.035 0.395 9.47 0.555 ;
      RECT 8.71 1.195 8.91 1.355 ;
      RECT 8.91 0.775 9.05 1.345 ;
      RECT 8.89 0.775 9.07 0.995 ;
      RECT 8.38 1.605 9.06 1.805 ;
      RECT 8.38 0.785 8.54 1.805 ;
      RECT 7.035 1.98 8.13 2.14 ;
      RECT 7.97 0.785 8.13 2.14 ;
      RECT 7.035 1.605 7.195 2.14 ;
      RECT 6.515 1.18 6.675 1.805 ;
      RECT 6.105 1.18 6.675 1.34 ;
      RECT 6.105 0.785 6.265 1.34 ;
      RECT 4.245 0.41 4.405 0.985 ;
      RECT 4.21 0.41 4.43 0.59 ;
      RECT 5.825 0.41 6.025 0.57 ;
      RECT 4.21 0.42 6.025 0.56 ;
      RECT 4.245 1.18 4.405 1.805 ;
      RECT 4.245 1.18 4.815 1.34 ;
      RECT 4.655 0.785 4.815 1.34 ;
      RECT 4.655 0.785 5.335 0.985 ;
      RECT 4.92 1.96 5.12 2.15 ;
      RECT 4.91 1.96 5.13 2.14 ;
      RECT 4.91 1.96 5.335 2.12 ;
      RECT 5.175 1.605 5.335 2.12 ;
      RECT 4.61 1.5 4.855 1.805 ;
      RECT 4.565 1.5 5.015 1.8 ;
      RECT 2.565 0.725 2.745 2.135 ;
      RECT 2.585 0.39 2.745 2.135 ;
      RECT 3.405 0.39 3.565 2.13 ;
      RECT 2.55 0.725 2.775 2.13 ;
      RECT 2.55 1.74 3.565 1.9 ;
      RECT 2.985 1.36 3.165 1.58 ;
      RECT 2.995 0.66 3.155 1.58 ;
      RECT 1.355 0.39 1.515 2.13 ;
      RECT 0.505 0.43 0.725 2.13 ;
      RECT 0.505 1.74 1.515 1.9 ;
      RECT 0.535 0.39 0.695 2.13 ;
      RECT 12.095 0.785 12.775 0.985 ;
      RECT 11.165 1.605 11.845 1.805 ;
      RECT 10.425 0.39 10.87 0.625 ;
      RECT 6.92 1.165 7.435 1.385 ;
      RECT 6.48 0.645 6.775 0.995 ;
      RECT 5.585 1.605 6.285 1.805 ;
      RECT 5.505 0.765 5.81 1.12 ;
    LAYER V12 ;
      RECT 13.035 0.815 13.175 0.955 ;
      RECT 12.375 1.99 12.515 2.13 ;
      RECT 10.51 0.44 10.65 0.58 ;
      RECT 9.605 1.99 9.745 2.13 ;
      RECT 8.91 0.815 9.05 0.955 ;
      RECT 7.255 1.21 7.395 1.35 ;
      RECT 6.525 0.815 6.665 0.955 ;
      RECT 5.595 0.815 5.735 0.955 ;
      RECT 4.95 1.98 5.09 2.12 ;
      RECT 4.665 1.635 4.805 1.775 ;
      RECT 4.25 0.43 4.39 0.57 ;
      RECT 3.005 1.4 3.145 1.54 ;
      RECT 2.595 1.045 2.735 1.185 ;
      RECT 2.595 1.35 2.735 1.49 ;
      RECT 2.59 0.745 2.73 0.885 ;
      RECT 2.59 1.675 2.73 1.815 ;
      RECT 2.585 1.955 2.725 2.095 ;
      RECT 0.545 0.45 0.685 0.59 ;
      RECT 0.545 0.73 0.685 0.87 ;
      RECT 0.545 1.4 0.685 1.54 ;
      RECT 0.545 1.69 0.685 1.83 ;
      RECT 0.545 1.97 0.685 2.11 ;
    LAYER M2 ;
      RECT 0.505 0.155 0.725 2.15 ;
      RECT 2.965 1.38 3.185 1.56 ;
      RECT 3.005 0.155 3.145 1.56 ;
      RECT 13.015 0.775 13.195 0.995 ;
      RECT 8.87 0.795 9.09 0.975 ;
      RECT 8.91 0.145 9.05 0.975 ;
      RECT 13.035 0.25 13.175 0.995 ;
      RECT 10.49 0.16 10.67 0.62 ;
      RECT 4.23 0.16 4.985 0.61 ;
      RECT 3.005 0.16 4.985 0.565 ;
      RECT 0.5 0.25 13.175 0.39 ;
      RECT 0.5 0.16 12.9 0.39 ;
      RECT 0.5 0.155 4.335 0.39 ;
      RECT 2.545 2.055 12.505 2.285 ;
      RECT 12.355 1.95 12.535 2.17 ;
      RECT 9.585 1.95 9.765 2.285 ;
      RECT 4.93 1.94 5.11 2.285 ;
      RECT 2.545 1.95 4.485 2.285 ;
      RECT 2.545 1.935 2.78 2.285 ;
      RECT 2.55 0.705 2.78 2.285 ;
      RECT 4.645 1.595 4.825 1.815 ;
      RECT 4.665 1.19 4.805 1.815 ;
      RECT 7.235 1.17 7.415 1.39 ;
      RECT 4.665 1.19 7.415 1.33 ;
      RECT 6.525 0.775 6.665 1.33 ;
      RECT 5.595 0.775 5.735 1.33 ;
      RECT 6.505 0.775 6.685 0.995 ;
      RECT 5.575 0.775 5.755 0.995 ;
  END
END dig_poly_XOR_BUF2_x1

END LIBRARY
