/*
:set expandtab
:set tabstop=4
:set shiftwidth=4
:retab

*/

`include "ahbl_defines.vh"

package ahbl_bus_mux_common;



endpackage : ahbl_bus_mux_common
