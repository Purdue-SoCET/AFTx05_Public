VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ring_161x
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ring_161x 0 0 ;
  SIZE 34.44 BY 15.36 ;
  SYMMETRY X Y ;
  SITE CoreSite8T ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 34.44 0.23 ;
        RECT 34.155 0 34.315 0.76 ;
        RECT 33.335 0 33.495 0.5 ;
        RECT 32.925 0 33.085 0.76 ;
        RECT 32.105 0 32.265 0.5 ;
        RECT 31.695 0 31.855 0.76 ;
        RECT 30.875 0 31.035 0.5 ;
        RECT 30.465 0 30.625 0.76 ;
        RECT 29.645 0 29.805 0.5 ;
        RECT 29.235 0 29.395 0.76 ;
        RECT 28.415 0 28.575 0.5 ;
        RECT 28.005 0 28.165 0.76 ;
        RECT 27.185 0 27.345 0.5 ;
        RECT 26.775 0 26.935 0.76 ;
        RECT 25.955 0 26.115 0.5 ;
        RECT 25.545 0 25.705 0.76 ;
        RECT 24.725 0 24.885 0.5 ;
        RECT 24.315 0 24.475 0.76 ;
        RECT 23.495 0 23.655 0.5 ;
        RECT 23.085 0 23.245 0.76 ;
        RECT 22.265 0 22.425 0.5 ;
        RECT 21.855 0 22.015 0.76 ;
        RECT 21.035 0 21.195 0.5 ;
        RECT 20.625 0 20.785 0.76 ;
        RECT 19.805 0 19.965 0.5 ;
        RECT 19.395 0 19.555 0.76 ;
        RECT 18.575 0 18.735 0.5 ;
        RECT 18.165 0 18.325 0.76 ;
        RECT 17.345 0 17.505 0.5 ;
        RECT 16.935 0 17.095 0.76 ;
        RECT 16.115 0 16.275 0.5 ;
        RECT 15.705 0 15.865 0.76 ;
        RECT 14.885 0 15.045 0.5 ;
        RECT 14.475 0 14.635 0.76 ;
        RECT 13.655 0 13.815 0.5 ;
        RECT 13.245 0 13.405 0.76 ;
        RECT 12.425 0 12.585 0.5 ;
        RECT 12.015 0 12.175 0.76 ;
        RECT 11.195 0 11.355 0.5 ;
        RECT 10.785 0 10.945 0.76 ;
        RECT 9.965 0 10.125 0.5 ;
        RECT 9.555 0 9.715 0.76 ;
        RECT 8.735 0 8.895 0.5 ;
        RECT 8.325 0 8.485 0.76 ;
        RECT 7.505 0 7.665 0.5 ;
        RECT 7.095 0 7.255 0.76 ;
        RECT 6.275 0 6.435 0.5 ;
        RECT 5.865 0 6.025 0.76 ;
        RECT 5.045 0 5.205 0.5 ;
        RECT 4.635 0 4.795 0.76 ;
        RECT 3.815 0 3.975 0.5 ;
        RECT 3.405 0 3.565 0.76 ;
        RECT 2.585 0 2.745 0.5 ;
        RECT 2.175 0 2.335 0.76 ;
        RECT 1.355 0 1.515 0.5 ;
        RECT 0.945 0 1.105 0.76 ;
        RECT 0 4.89 34.44 5.35 ;
        RECT 34.155 4.62 34.315 5.88 ;
        RECT 33.335 4.36 33.495 5.62 ;
        RECT 32.925 4.62 33.085 5.88 ;
        RECT 32.105 4.36 32.265 5.62 ;
        RECT 31.695 4.62 31.855 5.88 ;
        RECT 30.875 4.36 31.035 5.62 ;
        RECT 30.465 4.62 30.625 5.88 ;
        RECT 29.645 4.36 29.805 5.62 ;
        RECT 29.235 4.62 29.395 5.88 ;
        RECT 28.415 4.36 28.575 5.62 ;
        RECT 28.005 4.62 28.165 5.88 ;
        RECT 27.185 4.36 27.345 5.62 ;
        RECT 26.775 4.62 26.935 5.88 ;
        RECT 25.955 4.36 26.115 5.62 ;
        RECT 25.545 4.62 25.705 5.88 ;
        RECT 24.725 4.36 24.885 5.62 ;
        RECT 24.315 4.62 24.475 5.88 ;
        RECT 23.495 4.36 23.655 5.62 ;
        RECT 23.085 4.62 23.245 5.88 ;
        RECT 22.265 4.36 22.425 5.62 ;
        RECT 21.855 4.62 22.015 5.88 ;
        RECT 21.035 4.36 21.195 5.62 ;
        RECT 20.625 4.62 20.785 5.88 ;
        RECT 19.805 4.36 19.965 5.62 ;
        RECT 19.395 4.62 19.555 5.88 ;
        RECT 18.575 4.36 18.735 5.62 ;
        RECT 18.165 4.62 18.325 5.88 ;
        RECT 17.345 4.36 17.505 5.62 ;
        RECT 16.935 4.62 17.095 5.88 ;
        RECT 16.115 4.36 16.275 5.62 ;
        RECT 15.705 4.62 15.865 5.88 ;
        RECT 14.885 4.36 15.045 5.62 ;
        RECT 14.475 4.62 14.635 5.88 ;
        RECT 13.655 4.36 13.815 5.62 ;
        RECT 13.245 4.62 13.405 5.88 ;
        RECT 12.425 4.36 12.585 5.62 ;
        RECT 12.015 4.62 12.175 5.88 ;
        RECT 11.195 4.36 11.355 5.62 ;
        RECT 10.785 4.62 10.945 5.88 ;
        RECT 9.965 4.36 10.125 5.62 ;
        RECT 9.555 4.62 9.715 5.88 ;
        RECT 8.735 4.36 8.895 5.62 ;
        RECT 8.325 4.62 8.485 5.88 ;
        RECT 7.505 4.36 7.665 5.62 ;
        RECT 7.095 4.62 7.255 5.88 ;
        RECT 6.275 4.36 6.435 5.62 ;
        RECT 5.865 4.62 6.025 5.88 ;
        RECT 5.045 4.36 5.205 5.62 ;
        RECT 4.635 4.62 4.795 5.88 ;
        RECT 3.815 4.36 3.975 5.62 ;
        RECT 3.405 4.62 3.565 5.88 ;
        RECT 2.585 4.36 2.745 5.62 ;
        RECT 2.175 4.62 2.335 5.88 ;
        RECT 1.355 4.36 1.515 5.62 ;
        RECT 0.945 4.62 1.105 5.88 ;
        RECT 0.125 4.36 0.285 5.62 ;
        RECT 0 10.01 34.44 10.47 ;
        RECT 34.155 9.74 34.315 11 ;
        RECT 33.335 9.48 33.495 10.74 ;
        RECT 32.925 9.74 33.085 11 ;
        RECT 32.105 9.48 32.265 10.74 ;
        RECT 31.695 9.74 31.855 11 ;
        RECT 30.875 9.48 31.035 10.74 ;
        RECT 30.465 9.74 30.625 11 ;
        RECT 29.645 9.48 29.805 10.74 ;
        RECT 29.235 9.74 29.395 11 ;
        RECT 28.415 9.48 28.575 10.74 ;
        RECT 28.005 9.74 28.165 11 ;
        RECT 27.185 9.48 27.345 10.74 ;
        RECT 26.775 9.74 26.935 11 ;
        RECT 25.955 9.48 26.115 10.74 ;
        RECT 25.545 9.74 25.705 11 ;
        RECT 24.725 9.48 24.885 10.74 ;
        RECT 24.315 9.74 24.475 11 ;
        RECT 23.495 9.48 23.655 10.74 ;
        RECT 23.085 9.74 23.245 11 ;
        RECT 22.265 9.48 22.425 10.74 ;
        RECT 21.855 9.74 22.015 11 ;
        RECT 21.035 9.48 21.195 10.74 ;
        RECT 20.625 9.74 20.785 11 ;
        RECT 19.805 9.48 19.965 10.74 ;
        RECT 19.395 9.74 19.555 11 ;
        RECT 18.575 9.48 18.735 10.74 ;
        RECT 18.165 9.74 18.325 11 ;
        RECT 17.345 9.48 17.505 10.74 ;
        RECT 16.935 9.74 17.095 11 ;
        RECT 16.115 9.48 16.275 10.74 ;
        RECT 15.705 9.74 15.865 11 ;
        RECT 14.885 9.48 15.045 10.74 ;
        RECT 14.475 9.74 14.635 11 ;
        RECT 13.655 9.48 13.815 10.74 ;
        RECT 13.245 9.74 13.405 11 ;
        RECT 12.425 9.48 12.585 10.74 ;
        RECT 12.015 9.74 12.175 11 ;
        RECT 11.195 9.48 11.355 10.74 ;
        RECT 10.785 9.74 10.945 11 ;
        RECT 9.965 9.48 10.125 10.74 ;
        RECT 9.555 9.74 9.715 11 ;
        RECT 8.735 9.48 8.895 10.74 ;
        RECT 8.325 9.74 8.485 11 ;
        RECT 7.505 9.48 7.665 10.74 ;
        RECT 7.095 9.74 7.255 11 ;
        RECT 6.275 9.48 6.435 10.74 ;
        RECT 5.865 9.74 6.025 11 ;
        RECT 5.045 9.48 5.205 10.74 ;
        RECT 4.635 9.74 4.795 11 ;
        RECT 3.815 9.48 3.975 10.74 ;
        RECT 3.405 9.74 3.565 11 ;
        RECT 2.585 9.48 2.745 10.74 ;
        RECT 2.175 9.74 2.335 11 ;
        RECT 1.355 9.48 1.515 10.74 ;
        RECT 0.945 9.74 1.105 11 ;
        RECT 0.125 9.48 0.285 10.74 ;
        RECT 0 15.13 34.44 15.36 ;
        RECT 34.155 14.86 34.315 15.36 ;
        RECT 33.335 14.6 33.495 15.36 ;
        RECT 32.925 14.86 33.085 15.36 ;
        RECT 32.105 14.6 32.265 15.36 ;
        RECT 31.695 14.86 31.855 15.36 ;
        RECT 30.875 14.6 31.035 15.36 ;
        RECT 30.465 14.86 30.625 15.36 ;
        RECT 29.645 14.6 29.805 15.36 ;
        RECT 29.235 14.86 29.395 15.36 ;
        RECT 28.415 14.6 28.575 15.36 ;
        RECT 28.005 14.86 28.165 15.36 ;
        RECT 27.185 14.6 27.345 15.36 ;
        RECT 26.775 14.86 26.935 15.36 ;
        RECT 25.955 14.6 26.115 15.36 ;
        RECT 25.545 14.86 25.705 15.36 ;
        RECT 24.725 14.6 24.885 15.36 ;
        RECT 24.315 14.86 24.475 15.36 ;
        RECT 23.495 14.6 23.655 15.36 ;
        RECT 23.085 14.86 23.245 15.36 ;
        RECT 22.265 14.6 22.425 15.36 ;
        RECT 21.855 14.86 22.015 15.36 ;
        RECT 21.035 14.6 21.195 15.36 ;
        RECT 20.625 14.86 20.785 15.36 ;
        RECT 19.805 14.6 19.965 15.36 ;
        RECT 19.395 14.86 19.555 15.36 ;
        RECT 18.575 14.6 18.735 15.36 ;
        RECT 18.165 14.86 18.325 15.36 ;
        RECT 17.345 14.6 17.505 15.36 ;
        RECT 16.935 14.86 17.095 15.36 ;
        RECT 16.115 14.6 16.275 15.36 ;
        RECT 15.705 14.86 15.865 15.36 ;
        RECT 14.885 14.6 15.045 15.36 ;
        RECT 14.475 14.86 14.635 15.36 ;
        RECT 13.655 14.6 13.815 15.36 ;
        RECT 13.245 14.86 13.405 15.36 ;
        RECT 12.425 14.6 12.585 15.36 ;
        RECT 12.015 14.86 12.175 15.36 ;
        RECT 11.195 14.6 11.355 15.36 ;
        RECT 10.785 14.86 10.945 15.36 ;
        RECT 9.965 14.6 10.125 15.36 ;
        RECT 9.555 14.86 9.715 15.36 ;
        RECT 8.735 14.6 8.895 15.36 ;
        RECT 8.325 14.86 8.485 15.36 ;
        RECT 7.505 14.86 7.665 15.36 ;
        RECT 6.685 14.6 6.845 15.36 ;
        RECT 6.275 14.6 6.435 15.36 ;
        RECT 5.455 14.86 5.615 15.36 ;
        RECT 4.635 14.6 4.795 15.36 ;
        RECT 4.225 14.6 4.385 15.36 ;
        RECT 3.405 14.6 3.565 15.36 ;
        RECT 2.585 14.6 2.745 15.36 ;
        RECT 1.765 14.6 1.925 15.36 ;
        RECT 0.945 14.6 1.105 15.36 ;
      LAYER M2 ;
        RECT 2.46 5.12 3.575 5.35 ;
        RECT 2.46 10.24 3.575 10.47 ;
        RECT 0 0 1.115 0.23 ;
        RECT 0 15.13 1.115 15.36 ;
      LAYER M3 ;
        RECT 2.46 5.12 3.575 5.35 ;
        RECT 2.46 10.24 3.575 10.47 ;
        RECT 0 0 1.115 0.23 ;
        RECT 0 15.13 1.115 15.36 ;
      LAYER V12 ;
        RECT 0.075 15.17 0.215 15.31 ;
        RECT 0.075 0.04 0.215 0.18 ;
        RECT 0.355 15.17 0.495 15.31 ;
        RECT 0.355 0.04 0.495 0.18 ;
        RECT 0.635 15.17 0.775 15.31 ;
        RECT 0.635 0.04 0.775 0.18 ;
        RECT 0.915 15.17 1.055 15.31 ;
        RECT 0.915 0.04 1.055 0.18 ;
        RECT 2.535 10.28 2.675 10.42 ;
        RECT 2.535 5.16 2.675 5.3 ;
        RECT 2.815 10.28 2.955 10.42 ;
        RECT 2.815 5.16 2.955 5.3 ;
        RECT 3.095 10.28 3.235 10.42 ;
        RECT 3.095 5.16 3.235 5.3 ;
        RECT 3.375 10.28 3.515 10.42 ;
        RECT 3.375 5.16 3.515 5.3 ;
      LAYER V23 ;
        RECT 0.075 15.17 0.215 15.31 ;
        RECT 0.075 0.04 0.215 0.18 ;
        RECT 0.355 15.17 0.495 15.31 ;
        RECT 0.355 0.04 0.495 0.18 ;
        RECT 0.635 15.17 0.775 15.31 ;
        RECT 0.635 0.04 0.775 0.18 ;
        RECT 0.915 15.17 1.055 15.31 ;
        RECT 0.915 0.04 1.055 0.18 ;
        RECT 2.535 10.28 2.675 10.42 ;
        RECT 2.535 5.16 2.675 5.3 ;
        RECT 2.815 10.28 2.955 10.42 ;
        RECT 2.815 5.16 2.955 5.3 ;
        RECT 3.095 10.28 3.235 10.42 ;
        RECT 3.095 5.16 3.235 5.3 ;
        RECT 3.375 10.28 3.515 10.42 ;
        RECT 3.375 5.16 3.515 5.3 ;
    END
  END vss!
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.115 0.71 0.295 1.77 ;
        RECT 0.125 0.71 0.285 1.81 ;
      LAYER M2 ;
        RECT 0.095 0.73 0.315 1.75 ;
      LAYER M3 ;
        RECT 0.115 0.71 0.295 1.77 ;
      LAYER V12 ;
        RECT 0.135 1.59 0.275 1.73 ;
        RECT 0.135 1.31 0.275 1.45 ;
        RECT 0.135 1.03 0.275 1.17 ;
        RECT 0.135 0.75 0.275 0.89 ;
      LAYER V23 ;
        RECT 0.135 1.59 0.275 1.73 ;
        RECT 0.135 1.31 0.275 1.45 ;
        RECT 0.135 1.03 0.275 1.17 ;
        RECT 0.135 0.75 0.275 0.89 ;
    END
  END EN
  PIN OUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.805 13.49 3.985 13.71 ;
        RECT 3.815 13.23 3.975 14.97 ;
        RECT 2.985 13.49 3.165 13.71 ;
        RECT 2.995 13.23 3.155 14.97 ;
        RECT 2.165 13.49 2.345 13.71 ;
        RECT 2.175 13.23 2.335 14.97 ;
        RECT 1.345 13.49 1.525 13.71 ;
        RECT 1.355 13.23 1.515 14.97 ;
      LAYER M2 ;
        RECT 3.785 13.51 4.005 13.69 ;
        RECT 1.325 13.53 4.005 13.67 ;
        RECT 2.05 13.51 3.185 13.69 ;
        RECT 1.325 13.51 1.545 13.69 ;
      LAYER M3 ;
        RECT 2.07 13.49 3.09 13.71 ;
      LAYER V12 ;
        RECT 1.365 13.53 1.505 13.67 ;
        RECT 2.185 13.53 2.325 13.67 ;
        RECT 3.005 13.53 3.145 13.67 ;
        RECT 3.825 13.53 3.965 13.67 ;
      LAYER V23 ;
        RECT 2.09 13.53 2.23 13.67 ;
        RECT 2.37 13.53 2.51 13.67 ;
        RECT 2.65 13.53 2.79 13.67 ;
        RECT 2.93 13.53 3.07 13.67 ;
    END
  END OUT
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.33 34.44 2.79 ;
        RECT 34.155 1.54 34.315 3.06 ;
        RECT 33.335 2.06 33.495 3.58 ;
        RECT 32.925 1.54 33.085 3.06 ;
        RECT 32.105 2.06 32.265 3.58 ;
        RECT 31.695 1.54 31.855 3.06 ;
        RECT 30.875 2.06 31.035 3.58 ;
        RECT 30.465 1.54 30.625 3.06 ;
        RECT 29.645 2.06 29.805 3.58 ;
        RECT 29.235 1.54 29.395 3.06 ;
        RECT 28.415 2.06 28.575 3.58 ;
        RECT 28.005 1.54 28.165 3.06 ;
        RECT 27.185 2.06 27.345 3.58 ;
        RECT 26.775 1.54 26.935 3.06 ;
        RECT 25.955 2.06 26.115 3.58 ;
        RECT 25.545 1.54 25.705 3.06 ;
        RECT 24.725 2.06 24.885 3.58 ;
        RECT 24.315 1.54 24.475 3.06 ;
        RECT 23.495 2.06 23.655 3.58 ;
        RECT 23.085 1.54 23.245 3.06 ;
        RECT 22.265 2.06 22.425 3.58 ;
        RECT 21.855 1.54 22.015 3.06 ;
        RECT 21.035 2.06 21.195 3.58 ;
        RECT 20.625 1.54 20.785 3.06 ;
        RECT 19.805 2.06 19.965 3.58 ;
        RECT 19.395 1.54 19.555 3.06 ;
        RECT 18.575 2.06 18.735 3.58 ;
        RECT 18.165 1.54 18.325 3.06 ;
        RECT 17.345 2.06 17.505 3.58 ;
        RECT 16.935 1.54 17.095 3.06 ;
        RECT 16.115 2.06 16.275 3.58 ;
        RECT 15.705 1.54 15.865 3.06 ;
        RECT 14.885 2.06 15.045 3.58 ;
        RECT 14.475 1.54 14.635 3.06 ;
        RECT 13.655 2.06 13.815 3.58 ;
        RECT 13.245 1.54 13.405 3.06 ;
        RECT 12.425 2.06 12.585 3.58 ;
        RECT 12.015 1.54 12.175 3.06 ;
        RECT 11.195 2.06 11.355 3.58 ;
        RECT 10.785 1.54 10.945 3.06 ;
        RECT 9.965 2.06 10.125 3.58 ;
        RECT 9.555 1.54 9.715 3.06 ;
        RECT 8.735 2.06 8.895 3.58 ;
        RECT 8.325 1.54 8.485 3.06 ;
        RECT 7.505 2.06 7.665 3.58 ;
        RECT 7.095 1.54 7.255 3.06 ;
        RECT 6.275 2.06 6.435 3.58 ;
        RECT 5.865 1.54 6.025 3.06 ;
        RECT 5.045 2.06 5.205 3.58 ;
        RECT 4.635 1.54 4.795 3.06 ;
        RECT 3.815 2.06 3.975 3.58 ;
        RECT 3.405 1.54 3.565 3.06 ;
        RECT 2.585 2.06 2.745 3.58 ;
        RECT 2.175 1.54 2.335 3.06 ;
        RECT 1.355 2.06 1.515 3.58 ;
        RECT 0.945 1.97 1.105 3.06 ;
        RECT 0.125 1.97 0.285 3.58 ;
        RECT 0 7.45 34.44 7.91 ;
        RECT 34.155 6.66 34.315 8.18 ;
        RECT 33.335 7.18 33.495 8.7 ;
        RECT 32.925 6.66 33.085 8.18 ;
        RECT 32.105 7.18 32.265 8.7 ;
        RECT 31.695 6.66 31.855 8.18 ;
        RECT 30.875 7.18 31.035 8.7 ;
        RECT 30.465 6.66 30.625 8.18 ;
        RECT 29.645 7.18 29.805 8.7 ;
        RECT 29.235 6.66 29.395 8.18 ;
        RECT 28.415 7.18 28.575 8.7 ;
        RECT 28.005 6.66 28.165 8.18 ;
        RECT 27.185 7.18 27.345 8.7 ;
        RECT 26.775 6.66 26.935 8.18 ;
        RECT 25.955 7.18 26.115 8.7 ;
        RECT 25.545 6.66 25.705 8.18 ;
        RECT 24.725 7.18 24.885 8.7 ;
        RECT 24.315 6.66 24.475 8.18 ;
        RECT 23.495 7.18 23.655 8.7 ;
        RECT 23.085 6.66 23.245 8.18 ;
        RECT 22.265 7.18 22.425 8.7 ;
        RECT 21.855 6.66 22.015 8.18 ;
        RECT 21.035 7.18 21.195 8.7 ;
        RECT 20.625 6.66 20.785 8.18 ;
        RECT 19.805 7.18 19.965 8.7 ;
        RECT 19.395 6.66 19.555 8.18 ;
        RECT 18.575 7.18 18.735 8.7 ;
        RECT 18.165 6.66 18.325 8.18 ;
        RECT 17.345 7.18 17.505 8.7 ;
        RECT 16.935 6.66 17.095 8.18 ;
        RECT 16.115 7.18 16.275 8.7 ;
        RECT 15.705 6.66 15.865 8.18 ;
        RECT 14.885 7.18 15.045 8.7 ;
        RECT 14.475 6.66 14.635 8.18 ;
        RECT 13.655 7.18 13.815 8.7 ;
        RECT 13.245 6.66 13.405 8.18 ;
        RECT 12.425 7.18 12.585 8.7 ;
        RECT 12.015 6.66 12.175 8.18 ;
        RECT 11.195 7.18 11.355 8.7 ;
        RECT 10.785 6.66 10.945 8.18 ;
        RECT 9.965 7.18 10.125 8.7 ;
        RECT 9.555 6.66 9.715 8.18 ;
        RECT 8.735 7.18 8.895 8.7 ;
        RECT 8.325 6.66 8.485 8.18 ;
        RECT 7.505 7.18 7.665 8.7 ;
        RECT 7.095 6.66 7.255 8.18 ;
        RECT 6.275 7.18 6.435 8.7 ;
        RECT 5.865 6.66 6.025 8.18 ;
        RECT 5.045 7.18 5.205 8.7 ;
        RECT 4.635 6.66 4.795 8.18 ;
        RECT 3.815 7.18 3.975 8.7 ;
        RECT 3.405 6.66 3.565 8.18 ;
        RECT 2.585 7.18 2.745 8.7 ;
        RECT 2.175 6.66 2.335 8.18 ;
        RECT 1.355 7.18 1.515 8.7 ;
        RECT 0.945 6.66 1.105 8.18 ;
        RECT 0.125 7.18 0.285 8.7 ;
        RECT 0 12.57 34.44 13.03 ;
        RECT 34.155 11.78 34.315 13.3 ;
        RECT 33.335 12.3 33.495 13.82 ;
        RECT 32.925 11.78 33.085 13.3 ;
        RECT 32.105 12.3 32.265 13.82 ;
        RECT 31.695 11.78 31.855 13.3 ;
        RECT 30.875 12.3 31.035 13.82 ;
        RECT 30.465 11.78 30.625 13.3 ;
        RECT 29.645 12.3 29.805 13.82 ;
        RECT 29.235 11.78 29.395 13.3 ;
        RECT 28.415 12.3 28.575 13.82 ;
        RECT 28.005 11.78 28.165 13.3 ;
        RECT 27.185 12.3 27.345 13.82 ;
        RECT 26.775 11.78 26.935 13.3 ;
        RECT 25.955 12.3 26.115 13.82 ;
        RECT 25.545 11.78 25.705 13.3 ;
        RECT 24.725 12.3 24.885 13.82 ;
        RECT 24.315 11.78 24.475 13.3 ;
        RECT 23.495 12.3 23.655 13.82 ;
        RECT 23.085 11.78 23.245 13.3 ;
        RECT 22.265 12.3 22.425 13.82 ;
        RECT 21.855 11.78 22.015 13.3 ;
        RECT 21.035 12.3 21.195 13.82 ;
        RECT 20.625 11.78 20.785 13.3 ;
        RECT 19.805 12.3 19.965 13.82 ;
        RECT 19.395 11.78 19.555 13.3 ;
        RECT 18.575 12.3 18.735 13.82 ;
        RECT 18.165 11.78 18.325 13.3 ;
        RECT 17.345 12.3 17.505 13.82 ;
        RECT 16.935 11.78 17.095 13.3 ;
        RECT 16.115 12.3 16.275 13.82 ;
        RECT 15.705 11.78 15.865 13.3 ;
        RECT 14.885 12.3 15.045 13.82 ;
        RECT 14.475 11.78 14.635 13.3 ;
        RECT 13.655 12.3 13.815 13.82 ;
        RECT 13.245 11.78 13.405 13.3 ;
        RECT 12.425 12.3 12.585 13.82 ;
        RECT 12.015 11.78 12.175 13.3 ;
        RECT 11.195 12.3 11.355 13.82 ;
        RECT 10.785 11.78 10.945 13.3 ;
        RECT 9.965 12.3 10.125 13.82 ;
        RECT 9.555 11.78 9.715 13.3 ;
        RECT 8.735 12.3 8.895 13.82 ;
        RECT 8.325 11.78 8.485 13.3 ;
        RECT 7.505 12.3 7.665 13.3 ;
        RECT 7.095 11.78 7.255 13.03 ;
        RECT 6.685 12.57 6.845 13.82 ;
        RECT 6.275 12.3 6.435 13.82 ;
        RECT 5.865 11.78 6.025 13.03 ;
        RECT 5.455 12.57 5.615 13.3 ;
        RECT 5.045 12.3 5.205 13.03 ;
        RECT 4.635 11.78 4.795 13.82 ;
        RECT 4.225 12.57 4.385 13.82 ;
        RECT 3.815 12.3 3.975 13.03 ;
        RECT 3.405 11.78 3.565 13.82 ;
        RECT 2.585 12.3 2.745 13.82 ;
        RECT 2.175 11.78 2.335 13.03 ;
        RECT 1.765 12.57 1.925 13.82 ;
        RECT 1.355 12.3 1.515 13.03 ;
        RECT 0.945 11.78 1.105 13.82 ;
        RECT 0.125 12.3 0.285 13.03 ;
      LAYER M2 ;
        RECT 9.89 2.56 11.005 2.79 ;
        RECT 9.89 7.68 11.005 7.91 ;
        RECT 9.89 12.8 11.005 13.03 ;
      LAYER M3 ;
        RECT 9.89 2.56 11.005 2.79 ;
        RECT 9.89 7.68 11.005 7.91 ;
        RECT 9.89 12.8 11.005 13.03 ;
      LAYER V12 ;
        RECT 9.965 12.84 10.105 12.98 ;
        RECT 9.965 7.72 10.105 7.86 ;
        RECT 9.965 2.6 10.105 2.74 ;
        RECT 10.245 12.84 10.385 12.98 ;
        RECT 10.245 7.72 10.385 7.86 ;
        RECT 10.245 2.6 10.385 2.74 ;
        RECT 10.525 12.84 10.665 12.98 ;
        RECT 10.525 7.72 10.665 7.86 ;
        RECT 10.525 2.6 10.665 2.74 ;
        RECT 10.805 12.84 10.945 12.98 ;
        RECT 10.805 7.72 10.945 7.86 ;
        RECT 10.805 2.6 10.945 2.74 ;
      LAYER V23 ;
        RECT 9.965 12.84 10.105 12.98 ;
        RECT 9.965 7.72 10.105 7.86 ;
        RECT 9.965 2.6 10.105 2.74 ;
        RECT 10.245 12.84 10.385 12.98 ;
        RECT 10.245 7.72 10.385 7.86 ;
        RECT 10.245 2.6 10.385 2.74 ;
        RECT 10.525 12.84 10.665 12.98 ;
        RECT 10.525 7.72 10.665 7.86 ;
        RECT 10.525 2.6 10.665 2.74 ;
        RECT 10.805 12.84 10.945 12.98 ;
        RECT 10.805 7.72 10.945 7.86 ;
        RECT 10.805 2.6 10.945 2.74 ;
    END
  END vdd!
  OBS
    LAYER M1 ;
      RECT 34.065 3.22 34.225 4.46 ;
      RECT 34.065 3.41 34.245 3.63 ;
      RECT 34.065 8.34 34.225 9.58 ;
      RECT 34.065 8.525 34.245 8.745 ;
      RECT 34.065 13.46 34.225 14.7 ;
      RECT 34.065 13.675 34.245 13.895 ;
      RECT 33.745 0.39 33.905 2.13 ;
      RECT 33.745 0.935 33.925 1.155 ;
      RECT 33.745 5.51 33.905 7.25 ;
      RECT 33.745 6.05 33.925 6.27 ;
      RECT 33.745 10.63 33.905 12.37 ;
      RECT 33.745 11.22 33.925 11.44 ;
      RECT 33.745 2.99 33.905 4.73 ;
      RECT 32.835 3.22 32.995 4.46 ;
      RECT 32.835 3.745 33.905 3.905 ;
      RECT 33.745 8.11 33.905 9.85 ;
      RECT 32.835 8.34 32.995 9.58 ;
      RECT 32.835 8.875 33.905 9.035 ;
      RECT 33.745 13.23 33.905 14.97 ;
      RECT 32.835 13.46 32.995 14.7 ;
      RECT 32.835 13.995 33.905 14.155 ;
      RECT 32.515 0.39 32.675 2.13 ;
      RECT 33.425 0.66 33.585 1.9 ;
      RECT 32.515 0.925 33.585 1.085 ;
      RECT 32.515 5.51 32.675 7.25 ;
      RECT 33.425 5.78 33.585 7.02 ;
      RECT 32.515 6.065 33.585 6.225 ;
      RECT 32.515 10.63 32.675 12.37 ;
      RECT 33.425 10.9 33.585 12.14 ;
      RECT 32.515 11.175 33.585 11.335 ;
      RECT 32.515 2.99 32.675 4.73 ;
      RECT 31.605 3.22 31.765 4.46 ;
      RECT 31.605 3.745 32.675 3.905 ;
      RECT 32.515 8.11 32.675 9.85 ;
      RECT 31.605 8.34 31.765 9.58 ;
      RECT 31.605 8.875 32.675 9.035 ;
      RECT 32.515 13.23 32.675 14.97 ;
      RECT 31.605 13.46 31.765 14.7 ;
      RECT 31.605 13.995 32.675 14.155 ;
      RECT 31.285 0.39 31.445 2.13 ;
      RECT 32.195 0.66 32.355 1.9 ;
      RECT 31.285 0.925 32.355 1.085 ;
      RECT 31.285 5.51 31.445 7.25 ;
      RECT 32.195 5.78 32.355 7.02 ;
      RECT 31.285 6.065 32.355 6.225 ;
      RECT 31.285 10.63 31.445 12.37 ;
      RECT 32.195 10.9 32.355 12.14 ;
      RECT 31.285 11.175 32.355 11.335 ;
      RECT 31.285 2.99 31.445 4.73 ;
      RECT 30.375 3.22 30.535 4.46 ;
      RECT 30.375 3.745 31.445 3.905 ;
      RECT 31.285 8.11 31.445 9.85 ;
      RECT 30.375 8.34 30.535 9.58 ;
      RECT 30.375 8.875 31.445 9.035 ;
      RECT 31.285 13.23 31.445 14.97 ;
      RECT 30.375 13.46 30.535 14.7 ;
      RECT 30.375 13.995 31.445 14.155 ;
      RECT 30.055 0.39 30.215 2.13 ;
      RECT 30.965 0.66 31.125 1.9 ;
      RECT 30.055 0.925 31.125 1.085 ;
      RECT 30.055 5.51 30.215 7.25 ;
      RECT 30.965 5.78 31.125 7.02 ;
      RECT 30.055 6.065 31.125 6.225 ;
      RECT 30.055 10.63 30.215 12.37 ;
      RECT 30.965 10.9 31.125 12.14 ;
      RECT 30.055 11.175 31.125 11.335 ;
      RECT 30.055 2.99 30.215 4.73 ;
      RECT 29.145 3.22 29.305 4.46 ;
      RECT 29.145 3.745 30.215 3.905 ;
      RECT 30.055 8.11 30.215 9.85 ;
      RECT 29.145 8.34 29.305 9.58 ;
      RECT 29.145 8.875 30.215 9.035 ;
      RECT 30.055 13.23 30.215 14.97 ;
      RECT 29.145 13.46 29.305 14.7 ;
      RECT 29.145 13.995 30.215 14.155 ;
      RECT 28.825 0.39 28.985 2.13 ;
      RECT 29.735 0.66 29.895 1.9 ;
      RECT 28.825 0.925 29.895 1.085 ;
      RECT 28.825 5.51 28.985 7.25 ;
      RECT 29.735 5.78 29.895 7.02 ;
      RECT 28.825 6.065 29.895 6.225 ;
      RECT 28.825 10.63 28.985 12.37 ;
      RECT 29.735 10.9 29.895 12.14 ;
      RECT 28.825 11.175 29.895 11.335 ;
      RECT 28.825 2.99 28.985 4.73 ;
      RECT 27.915 3.22 28.075 4.46 ;
      RECT 27.915 3.745 28.985 3.905 ;
      RECT 28.825 8.11 28.985 9.85 ;
      RECT 27.915 8.34 28.075 9.58 ;
      RECT 27.915 8.875 28.985 9.035 ;
      RECT 28.825 13.23 28.985 14.97 ;
      RECT 27.915 13.46 28.075 14.7 ;
      RECT 27.915 13.995 28.985 14.155 ;
      RECT 27.595 0.39 27.755 2.13 ;
      RECT 28.505 0.66 28.665 1.9 ;
      RECT 27.595 0.925 28.665 1.085 ;
      RECT 27.595 5.51 27.755 7.25 ;
      RECT 28.505 5.78 28.665 7.02 ;
      RECT 27.595 6.065 28.665 6.225 ;
      RECT 27.595 10.63 27.755 12.37 ;
      RECT 28.505 10.9 28.665 12.14 ;
      RECT 27.595 11.175 28.665 11.335 ;
      RECT 27.595 2.99 27.755 4.73 ;
      RECT 26.685 3.22 26.845 4.46 ;
      RECT 26.685 3.745 27.755 3.905 ;
      RECT 27.595 8.11 27.755 9.85 ;
      RECT 26.685 8.34 26.845 9.58 ;
      RECT 26.685 8.875 27.755 9.035 ;
      RECT 27.595 13.23 27.755 14.97 ;
      RECT 26.685 13.46 26.845 14.7 ;
      RECT 26.685 13.995 27.755 14.155 ;
      RECT 26.365 0.39 26.525 2.13 ;
      RECT 27.275 0.66 27.435 1.9 ;
      RECT 26.365 0.925 27.435 1.085 ;
      RECT 26.365 5.51 26.525 7.25 ;
      RECT 27.275 5.78 27.435 7.02 ;
      RECT 26.365 6.065 27.435 6.225 ;
      RECT 26.365 10.63 26.525 12.37 ;
      RECT 27.275 10.9 27.435 12.14 ;
      RECT 26.365 11.175 27.435 11.335 ;
      RECT 26.365 2.99 26.525 4.73 ;
      RECT 25.455 3.22 25.615 4.46 ;
      RECT 25.455 3.745 26.525 3.905 ;
      RECT 26.365 8.11 26.525 9.85 ;
      RECT 25.455 8.34 25.615 9.58 ;
      RECT 25.455 8.875 26.525 9.035 ;
      RECT 26.365 13.23 26.525 14.97 ;
      RECT 25.455 13.46 25.615 14.7 ;
      RECT 25.455 13.995 26.525 14.155 ;
      RECT 25.135 0.39 25.295 2.13 ;
      RECT 26.045 0.66 26.205 1.9 ;
      RECT 25.135 0.925 26.205 1.085 ;
      RECT 25.135 5.51 25.295 7.25 ;
      RECT 26.045 5.78 26.205 7.02 ;
      RECT 25.135 6.065 26.205 6.225 ;
      RECT 25.135 10.63 25.295 12.37 ;
      RECT 26.045 10.9 26.205 12.14 ;
      RECT 25.135 11.175 26.205 11.335 ;
      RECT 25.135 2.99 25.295 4.73 ;
      RECT 24.225 3.22 24.385 4.46 ;
      RECT 24.225 3.745 25.295 3.905 ;
      RECT 25.135 8.11 25.295 9.85 ;
      RECT 24.225 8.34 24.385 9.58 ;
      RECT 24.225 8.875 25.295 9.035 ;
      RECT 25.135 13.23 25.295 14.97 ;
      RECT 24.225 13.46 24.385 14.7 ;
      RECT 24.225 13.995 25.295 14.155 ;
      RECT 23.905 0.39 24.065 2.13 ;
      RECT 24.815 0.66 24.975 1.9 ;
      RECT 23.905 0.925 24.975 1.085 ;
      RECT 23.905 5.51 24.065 7.25 ;
      RECT 24.815 5.78 24.975 7.02 ;
      RECT 23.905 6.065 24.975 6.225 ;
      RECT 23.905 10.63 24.065 12.37 ;
      RECT 24.815 10.9 24.975 12.14 ;
      RECT 23.905 11.175 24.975 11.335 ;
      RECT 23.905 2.99 24.065 4.73 ;
      RECT 22.995 3.22 23.155 4.46 ;
      RECT 22.995 3.745 24.065 3.905 ;
      RECT 23.905 8.11 24.065 9.85 ;
      RECT 22.995 8.34 23.155 9.58 ;
      RECT 22.995 8.875 24.065 9.035 ;
      RECT 23.905 13.23 24.065 14.97 ;
      RECT 22.995 13.46 23.155 14.7 ;
      RECT 22.995 13.995 24.065 14.155 ;
      RECT 22.675 0.39 22.835 2.13 ;
      RECT 23.585 0.66 23.745 1.9 ;
      RECT 22.675 0.925 23.745 1.085 ;
      RECT 22.675 5.51 22.835 7.25 ;
      RECT 23.585 5.78 23.745 7.02 ;
      RECT 22.675 6.065 23.745 6.225 ;
      RECT 22.675 10.63 22.835 12.37 ;
      RECT 23.585 10.9 23.745 12.14 ;
      RECT 22.675 11.175 23.745 11.335 ;
      RECT 22.675 2.99 22.835 4.73 ;
      RECT 21.765 3.22 21.925 4.46 ;
      RECT 21.765 3.745 22.835 3.905 ;
      RECT 22.675 8.11 22.835 9.85 ;
      RECT 21.765 8.34 21.925 9.58 ;
      RECT 21.765 8.875 22.835 9.035 ;
      RECT 22.675 13.23 22.835 14.97 ;
      RECT 21.765 13.46 21.925 14.7 ;
      RECT 21.765 13.995 22.835 14.155 ;
      RECT 21.445 0.39 21.605 2.13 ;
      RECT 22.355 0.66 22.515 1.9 ;
      RECT 21.445 0.925 22.515 1.085 ;
      RECT 21.445 5.51 21.605 7.25 ;
      RECT 22.355 5.78 22.515 7.02 ;
      RECT 21.445 6.065 22.515 6.225 ;
      RECT 21.445 10.63 21.605 12.37 ;
      RECT 22.355 10.9 22.515 12.14 ;
      RECT 21.445 11.175 22.515 11.335 ;
      RECT 21.445 2.99 21.605 4.73 ;
      RECT 20.535 3.22 20.695 4.46 ;
      RECT 20.535 3.745 21.605 3.905 ;
      RECT 21.445 8.11 21.605 9.85 ;
      RECT 20.535 8.34 20.695 9.58 ;
      RECT 20.535 8.875 21.605 9.035 ;
      RECT 21.445 13.23 21.605 14.97 ;
      RECT 20.535 13.46 20.695 14.7 ;
      RECT 20.535 13.995 21.605 14.155 ;
      RECT 20.215 0.39 20.375 2.13 ;
      RECT 21.125 0.66 21.285 1.9 ;
      RECT 20.215 0.925 21.285 1.085 ;
      RECT 20.215 5.51 20.375 7.25 ;
      RECT 21.125 5.78 21.285 7.02 ;
      RECT 20.215 6.065 21.285 6.225 ;
      RECT 20.215 10.63 20.375 12.37 ;
      RECT 21.125 10.9 21.285 12.14 ;
      RECT 20.215 11.175 21.285 11.335 ;
      RECT 20.215 2.99 20.375 4.73 ;
      RECT 19.305 3.22 19.465 4.46 ;
      RECT 19.305 3.745 20.375 3.905 ;
      RECT 20.215 8.11 20.375 9.85 ;
      RECT 19.305 8.34 19.465 9.58 ;
      RECT 19.305 8.875 20.375 9.035 ;
      RECT 20.215 13.23 20.375 14.97 ;
      RECT 19.305 13.46 19.465 14.7 ;
      RECT 19.305 13.995 20.375 14.155 ;
      RECT 18.985 0.39 19.145 2.13 ;
      RECT 19.895 0.66 20.055 1.9 ;
      RECT 18.985 0.925 20.055 1.085 ;
      RECT 18.985 5.51 19.145 7.25 ;
      RECT 19.895 5.78 20.055 7.02 ;
      RECT 18.985 6.065 20.055 6.225 ;
      RECT 18.985 10.63 19.145 12.37 ;
      RECT 19.895 10.9 20.055 12.14 ;
      RECT 18.985 11.175 20.055 11.335 ;
      RECT 18.985 2.99 19.145 4.73 ;
      RECT 18.075 3.22 18.235 4.46 ;
      RECT 18.075 3.745 19.145 3.905 ;
      RECT 18.985 8.11 19.145 9.85 ;
      RECT 18.075 8.34 18.235 9.58 ;
      RECT 18.075 8.875 19.145 9.035 ;
      RECT 18.985 13.23 19.145 14.97 ;
      RECT 18.075 13.46 18.235 14.7 ;
      RECT 18.075 13.995 19.145 14.155 ;
      RECT 17.755 0.39 17.915 2.13 ;
      RECT 18.665 0.66 18.825 1.9 ;
      RECT 17.755 0.925 18.825 1.085 ;
      RECT 17.755 5.51 17.915 7.25 ;
      RECT 18.665 5.78 18.825 7.02 ;
      RECT 17.755 6.065 18.825 6.225 ;
      RECT 17.755 10.63 17.915 12.37 ;
      RECT 18.665 10.9 18.825 12.14 ;
      RECT 17.755 11.175 18.825 11.335 ;
      RECT 17.755 2.99 17.915 4.73 ;
      RECT 16.845 3.22 17.005 4.46 ;
      RECT 16.845 3.745 17.915 3.905 ;
      RECT 17.755 8.11 17.915 9.85 ;
      RECT 16.845 8.34 17.005 9.58 ;
      RECT 16.845 8.875 17.915 9.035 ;
      RECT 17.755 13.23 17.915 14.97 ;
      RECT 16.845 13.46 17.005 14.7 ;
      RECT 16.845 13.995 17.915 14.155 ;
      RECT 16.525 0.39 16.685 2.13 ;
      RECT 17.435 0.66 17.595 1.9 ;
      RECT 16.525 0.925 17.595 1.085 ;
      RECT 16.525 5.51 16.685 7.25 ;
      RECT 17.435 5.78 17.595 7.02 ;
      RECT 16.525 6.065 17.595 6.225 ;
      RECT 16.525 10.63 16.685 12.37 ;
      RECT 17.435 10.9 17.595 12.14 ;
      RECT 16.525 11.175 17.595 11.335 ;
      RECT 16.525 2.99 16.685 4.73 ;
      RECT 15.615 3.22 15.775 4.46 ;
      RECT 15.615 3.745 16.685 3.905 ;
      RECT 16.525 8.11 16.685 9.85 ;
      RECT 15.615 8.34 15.775 9.58 ;
      RECT 15.615 8.875 16.685 9.035 ;
      RECT 16.525 13.23 16.685 14.97 ;
      RECT 15.615 13.46 15.775 14.7 ;
      RECT 15.615 13.995 16.685 14.155 ;
      RECT 15.295 0.39 15.455 2.13 ;
      RECT 16.205 0.66 16.365 1.9 ;
      RECT 15.295 0.925 16.365 1.085 ;
      RECT 15.295 5.51 15.455 7.25 ;
      RECT 16.205 5.78 16.365 7.02 ;
      RECT 15.295 6.065 16.365 6.225 ;
      RECT 15.295 10.63 15.455 12.37 ;
      RECT 16.205 10.9 16.365 12.14 ;
      RECT 15.295 11.175 16.365 11.335 ;
      RECT 15.295 2.99 15.455 4.73 ;
      RECT 14.385 3.22 14.545 4.46 ;
      RECT 14.385 3.745 15.455 3.905 ;
      RECT 15.295 8.11 15.455 9.85 ;
      RECT 14.385 8.34 14.545 9.58 ;
      RECT 14.385 8.875 15.455 9.035 ;
      RECT 15.295 13.23 15.455 14.97 ;
      RECT 14.385 13.46 14.545 14.7 ;
      RECT 14.385 13.995 15.455 14.155 ;
      RECT 14.065 0.39 14.225 2.13 ;
      RECT 14.975 0.66 15.135 1.9 ;
      RECT 14.065 0.925 15.135 1.085 ;
      RECT 14.065 5.51 14.225 7.25 ;
      RECT 14.975 5.78 15.135 7.02 ;
      RECT 14.065 6.065 15.135 6.225 ;
      RECT 14.065 10.63 14.225 12.37 ;
      RECT 14.975 10.9 15.135 12.14 ;
      RECT 14.065 11.175 15.135 11.335 ;
      RECT 14.065 2.99 14.225 4.73 ;
      RECT 13.155 3.22 13.315 4.46 ;
      RECT 13.155 3.745 14.225 3.905 ;
      RECT 14.065 8.11 14.225 9.85 ;
      RECT 13.155 8.34 13.315 9.58 ;
      RECT 13.155 8.875 14.225 9.035 ;
      RECT 14.065 13.23 14.225 14.97 ;
      RECT 13.155 13.46 13.315 14.7 ;
      RECT 13.155 13.995 14.225 14.155 ;
      RECT 12.835 0.39 12.995 2.13 ;
      RECT 13.745 0.66 13.905 1.9 ;
      RECT 12.835 0.925 13.905 1.085 ;
      RECT 12.835 5.51 12.995 7.25 ;
      RECT 13.745 5.78 13.905 7.02 ;
      RECT 12.835 6.065 13.905 6.225 ;
      RECT 12.835 10.63 12.995 12.37 ;
      RECT 13.745 10.9 13.905 12.14 ;
      RECT 12.835 11.175 13.905 11.335 ;
      RECT 12.835 2.99 12.995 4.73 ;
      RECT 11.925 3.22 12.085 4.46 ;
      RECT 11.925 3.745 12.995 3.905 ;
      RECT 12.835 8.11 12.995 9.85 ;
      RECT 11.925 8.34 12.085 9.58 ;
      RECT 11.925 8.875 12.995 9.035 ;
      RECT 12.835 13.23 12.995 14.97 ;
      RECT 11.925 13.46 12.085 14.7 ;
      RECT 11.925 13.995 12.995 14.155 ;
      RECT 11.605 0.39 11.765 2.13 ;
      RECT 12.515 0.66 12.675 1.9 ;
      RECT 11.605 0.925 12.675 1.085 ;
      RECT 11.605 5.51 11.765 7.25 ;
      RECT 12.515 5.78 12.675 7.02 ;
      RECT 11.605 6.065 12.675 6.225 ;
      RECT 11.605 10.63 11.765 12.37 ;
      RECT 12.515 10.9 12.675 12.14 ;
      RECT 11.605 11.175 12.675 11.335 ;
      RECT 11.605 2.99 11.765 4.73 ;
      RECT 10.695 3.22 10.855 4.46 ;
      RECT 10.695 3.745 11.765 3.905 ;
      RECT 11.605 8.11 11.765 9.85 ;
      RECT 10.695 8.34 10.855 9.58 ;
      RECT 10.695 8.875 11.765 9.035 ;
      RECT 11.605 13.23 11.765 14.97 ;
      RECT 10.695 13.46 10.855 14.7 ;
      RECT 10.695 13.995 11.765 14.155 ;
      RECT 10.375 0.39 10.535 2.13 ;
      RECT 11.285 0.66 11.445 1.9 ;
      RECT 10.375 0.925 11.445 1.085 ;
      RECT 10.375 5.51 10.535 7.25 ;
      RECT 11.285 5.78 11.445 7.02 ;
      RECT 10.375 6.065 11.445 6.225 ;
      RECT 10.375 10.63 10.535 12.37 ;
      RECT 11.285 10.9 11.445 12.14 ;
      RECT 10.375 11.175 11.445 11.335 ;
      RECT 10.375 2.99 10.535 4.73 ;
      RECT 9.465 3.22 9.625 4.46 ;
      RECT 9.465 3.745 10.535 3.905 ;
      RECT 10.375 8.11 10.535 9.85 ;
      RECT 9.465 8.34 9.625 9.58 ;
      RECT 9.465 8.875 10.535 9.035 ;
      RECT 10.375 13.23 10.535 14.97 ;
      RECT 9.465 13.46 9.625 14.7 ;
      RECT 9.465 13.995 10.535 14.155 ;
      RECT 9.145 0.39 9.305 2.13 ;
      RECT 10.055 0.66 10.215 1.9 ;
      RECT 9.145 0.925 10.215 1.085 ;
      RECT 9.145 5.51 9.305 7.25 ;
      RECT 10.055 5.78 10.215 7.02 ;
      RECT 9.145 6.065 10.215 6.225 ;
      RECT 9.145 10.63 9.305 12.37 ;
      RECT 10.055 10.9 10.215 12.14 ;
      RECT 9.145 11.175 10.215 11.335 ;
      RECT 9.145 2.99 9.305 4.73 ;
      RECT 8.235 3.22 8.395 4.46 ;
      RECT 8.235 3.745 9.305 3.905 ;
      RECT 9.145 8.11 9.305 9.85 ;
      RECT 8.235 8.34 8.395 9.58 ;
      RECT 8.235 8.875 9.305 9.035 ;
      RECT 9.145 13.23 9.305 14.97 ;
      RECT 8.235 13.46 8.395 14.7 ;
      RECT 8.235 13.995 9.305 14.155 ;
      RECT 9.125 13.43 9.305 13.65 ;
      RECT 7.915 0.39 8.075 2.13 ;
      RECT 8.825 0.66 8.985 1.9 ;
      RECT 7.915 0.925 8.985 1.085 ;
      RECT 7.915 5.51 8.075 7.25 ;
      RECT 8.825 5.78 8.985 7.02 ;
      RECT 7.915 6.065 8.985 6.225 ;
      RECT 7.915 10.63 8.075 12.37 ;
      RECT 8.825 10.9 8.985 12.14 ;
      RECT 7.915 11.175 8.985 11.335 ;
      RECT 7.915 2.99 8.075 4.73 ;
      RECT 7.005 3.22 7.165 4.46 ;
      RECT 7.005 3.745 8.075 3.905 ;
      RECT 7.915 8.11 8.075 9.85 ;
      RECT 7.005 8.34 7.165 9.58 ;
      RECT 7.005 8.875 8.075 9.035 ;
      RECT 7.915 13.23 8.075 14.97 ;
      RECT 7.415 13.46 7.575 14.7 ;
      RECT 7.415 13.995 8.075 14.155 ;
      RECT 6.685 0.39 6.845 2.13 ;
      RECT 7.595 0.66 7.755 1.9 ;
      RECT 6.685 0.925 7.755 1.085 ;
      RECT 6.685 5.51 6.845 7.25 ;
      RECT 7.595 5.78 7.755 7.02 ;
      RECT 6.685 6.065 7.755 6.225 ;
      RECT 6.685 10.63 6.845 12.37 ;
      RECT 7.595 10.9 7.755 12.14 ;
      RECT 6.685 11.175 7.755 11.335 ;
      RECT 7.095 13.23 7.255 14.97 ;
      RECT 7.075 14.005 7.255 14.225 ;
      RECT 6.685 2.99 6.845 4.73 ;
      RECT 5.775 3.22 5.935 4.46 ;
      RECT 5.775 3.745 6.845 3.905 ;
      RECT 6.685 8.11 6.845 9.85 ;
      RECT 5.775 8.34 5.935 9.58 ;
      RECT 5.775 8.875 6.845 9.035 ;
      RECT 5.455 0.39 5.615 2.13 ;
      RECT 6.365 0.66 6.525 1.9 ;
      RECT 5.455 0.925 6.525 1.085 ;
      RECT 5.455 5.51 5.615 7.25 ;
      RECT 6.365 5.78 6.525 7.02 ;
      RECT 5.455 6.065 6.525 6.225 ;
      RECT 5.455 10.63 5.615 12.37 ;
      RECT 6.365 10.9 6.525 12.14 ;
      RECT 5.455 11.175 6.525 11.335 ;
      RECT 5.865 13.23 6.025 14.97 ;
      RECT 5.045 13.23 5.205 14.97 ;
      RECT 5.02 14.155 5.24 14.335 ;
      RECT 5.045 13.46 6.025 13.62 ;
      RECT 5.455 13.78 5.615 14.7 ;
      RECT 5.445 14.005 5.625 14.225 ;
      RECT 5.455 2.99 5.615 4.73 ;
      RECT 4.545 3.22 4.705 4.46 ;
      RECT 4.545 3.745 5.615 3.905 ;
      RECT 5.455 8.11 5.615 9.85 ;
      RECT 4.545 8.34 4.705 9.58 ;
      RECT 4.545 8.875 5.615 9.035 ;
      RECT 4.225 0.39 4.385 2.13 ;
      RECT 5.135 0.66 5.295 1.9 ;
      RECT 4.225 0.925 5.295 1.085 ;
      RECT 4.225 5.51 4.385 7.25 ;
      RECT 5.135 5.78 5.295 7.02 ;
      RECT 4.225 6.065 5.295 6.225 ;
      RECT 4.225 10.63 4.385 12.37 ;
      RECT 5.135 10.9 5.295 12.14 ;
      RECT 4.225 11.175 5.295 11.335 ;
      RECT 4.225 2.99 4.385 4.73 ;
      RECT 3.315 3.22 3.475 4.46 ;
      RECT 3.315 3.745 4.385 3.905 ;
      RECT 4.225 8.11 4.385 9.85 ;
      RECT 3.315 8.34 3.475 9.58 ;
      RECT 3.315 8.875 4.385 9.035 ;
      RECT 2.995 0.39 3.155 2.13 ;
      RECT 3.905 0.66 4.065 1.9 ;
      RECT 2.995 0.925 4.065 1.085 ;
      RECT 2.995 5.51 3.155 7.25 ;
      RECT 3.905 5.78 4.065 7.02 ;
      RECT 2.995 6.065 4.065 6.225 ;
      RECT 2.995 10.63 3.155 12.37 ;
      RECT 3.905 10.9 4.065 12.14 ;
      RECT 2.995 11.175 4.065 11.335 ;
      RECT 2.995 2.99 3.155 4.73 ;
      RECT 2.085 3.22 2.245 4.46 ;
      RECT 2.085 3.745 3.155 3.905 ;
      RECT 2.995 8.11 3.155 9.85 ;
      RECT 2.085 8.34 2.245 9.58 ;
      RECT 2.085 8.875 3.155 9.035 ;
      RECT 1.765 0.39 1.925 2.13 ;
      RECT 2.675 0.66 2.835 1.9 ;
      RECT 1.765 0.925 2.835 1.085 ;
      RECT 1.765 5.51 1.925 7.25 ;
      RECT 2.675 5.78 2.835 7.02 ;
      RECT 1.765 6.065 2.835 6.225 ;
      RECT 1.765 10.63 1.925 12.37 ;
      RECT 2.675 10.9 2.835 12.14 ;
      RECT 1.765 11.175 2.835 11.335 ;
      RECT 1.765 2.99 1.925 4.73 ;
      RECT 0.855 3.22 1.015 4.46 ;
      RECT 0.855 3.745 1.925 3.905 ;
      RECT 1.765 8.11 1.925 9.85 ;
      RECT 0.855 8.34 1.015 9.58 ;
      RECT 0.855 8.875 1.925 9.035 ;
      RECT 1.445 0.66 1.605 1.9 ;
      RECT 1.425 0.72 1.605 0.94 ;
      RECT 0.535 5.51 0.695 7.25 ;
      RECT 1.445 5.78 1.605 7.02 ;
      RECT 0.535 6.065 1.605 6.225 ;
      RECT 0.535 10.63 0.695 12.37 ;
      RECT 1.445 10.9 1.605 12.14 ;
      RECT 0.535 11.175 1.605 11.335 ;
      RECT 0.945 0.92 1.105 1.81 ;
      RECT 0.915 1.115 1.135 1.295 ;
      RECT 0.535 0.39 0.695 2.17 ;
      RECT 0.525 0.72 0.705 0.94 ;
      RECT 0.105 0.39 0.695 0.55 ;
      RECT 0.535 2.99 0.695 4.73 ;
      RECT 0.515 3.69 0.695 3.91 ;
      RECT 0.535 8.11 0.695 9.85 ;
      RECT 0.515 8.845 0.695 9.065 ;
      RECT 0.215 5.78 0.375 7.02 ;
      RECT 0.195 6.015 0.375 6.235 ;
      RECT 0.215 10.9 0.375 12.14 ;
      RECT 0.195 11.17 0.375 11.39 ;
      RECT 3.345 13.98 3.625 14.44 ;
      RECT 2.525 13.98 2.805 14.44 ;
      RECT 1.705 13.98 1.985 14.44 ;
    LAYER V12 ;
      RECT 34.085 3.45 34.225 3.59 ;
      RECT 34.085 8.565 34.225 8.705 ;
      RECT 34.085 13.715 34.225 13.855 ;
      RECT 33.765 0.975 33.905 1.115 ;
      RECT 33.765 6.09 33.905 6.23 ;
      RECT 33.765 11.26 33.905 11.4 ;
      RECT 9.145 13.47 9.285 13.61 ;
      RECT 7.095 14.045 7.235 14.185 ;
      RECT 5.465 14.045 5.605 14.185 ;
      RECT 5.06 14.175 5.2 14.315 ;
      RECT 3.415 14.17 3.555 14.31 ;
      RECT 2.595 14.17 2.735 14.31 ;
      RECT 1.775 14.17 1.915 14.31 ;
      RECT 1.445 0.76 1.585 0.9 ;
      RECT 0.955 1.135 1.095 1.275 ;
      RECT 0.545 0.76 0.685 0.9 ;
      RECT 0.535 3.73 0.675 3.87 ;
      RECT 0.535 8.885 0.675 9.025 ;
      RECT 0.215 6.055 0.355 6.195 ;
      RECT 0.215 11.21 0.355 11.35 ;
    LAYER M2 ;
      RECT 34.045 3.43 34.265 3.61 ;
      RECT 34.075 0.995 34.215 3.61 ;
      RECT 33.725 0.995 34.215 1.135 ;
      RECT 33.725 0.955 33.945 1.135 ;
      RECT 34.045 8.545 34.265 8.725 ;
      RECT 34.075 6.11 34.215 8.725 ;
      RECT 33.725 6.11 34.215 6.25 ;
      RECT 33.725 6.07 33.945 6.25 ;
      RECT 34.045 13.695 34.265 13.875 ;
      RECT 34.105 11.26 34.245 13.875 ;
      RECT 33.725 11.24 33.945 11.42 ;
      RECT 33.725 11.26 34.245 11.4 ;
      RECT 9.105 13.45 9.325 13.63 ;
      RECT 9.105 13.135 9.245 13.63 ;
      RECT 0.955 13.135 9.245 13.275 ;
      RECT 0.955 1.095 1.095 13.275 ;
      RECT 0.935 1.095 1.115 1.315 ;
      RECT 7.055 14.025 7.275 14.205 ;
      RECT 5.425 14.025 5.645 14.205 ;
      RECT 5.425 14.045 7.275 14.185 ;
      RECT 5.04 14.135 5.22 14.355 ;
      RECT 3.375 14.15 3.595 14.33 ;
      RECT 2.555 14.15 2.775 14.33 ;
      RECT 1.735 14.15 1.955 14.33 ;
      RECT 1.735 14.17 5.22 14.31 ;
      RECT 1.405 0.74 1.625 0.92 ;
      RECT 0.505 0.74 0.725 0.92 ;
      RECT 0.505 0.76 1.625 0.9 ;
      RECT 0.175 6.035 0.395 6.215 ;
      RECT 0.23 6.025 0.395 6.215 ;
      RECT 0.23 3.75 0.37 6.215 ;
      RECT 0.23 3.75 0.715 3.89 ;
      RECT 0.495 3.71 0.715 3.89 ;
      RECT 0.175 11.19 0.395 11.37 ;
      RECT 0.23 11.18 0.395 11.37 ;
      RECT 0.23 8.905 0.37 11.37 ;
      RECT 0.23 8.905 0.715 9.045 ;
      RECT 0.495 8.865 0.715 9.045 ;
  END
END ring_161x

END LIBRARY
